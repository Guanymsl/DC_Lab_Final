module bullet1_palette(output reg [23:0] color_map [0:15]);
    initial begin
        color_map[0] = 24'h000000; // Transparent
        color_map[1] = 24'hffffff;
        color_map[2] = 24'h7fffff;
        color_map[3] = 24'h8dfe8d;
        color_map[4] = 24'h77dbbd;
        color_map[5] = 24'h00ffff;
        color_map[6] = 24'h72ccbb;
        color_map[7] = 24'h71c6c2;
        color_map[8] = 24'h75c1c3;
        color_map[9] = 24'h72c0c8;
        color_map[10] = 24'h64c3bc;
        color_map[11] = 24'h5ebec0;
        color_map[12] = 24'h4db9be;
        color_map[13] = 24'h57aca9;
        color_map[14] = 24'h7f7f7f;
        color_map[15] = 24'h000000;
    end
endmodule

module bullet1_lut(output reg [3:0] pixel_data [0:24][0:24]);
    initial begin
        pixel_data[0][0] = 0;
        pixel_data[0][1] = 0;
        pixel_data[0][2] = 0;
        pixel_data[0][3] = 0;
        pixel_data[0][4] = 0;
        pixel_data[0][5] = 0;
        pixel_data[0][6] = 0;
        pixel_data[0][7] = 0;
        pixel_data[0][8] = 0;
        pixel_data[0][9] = 0;
        pixel_data[0][10] = 0;
        pixel_data[0][11] = 0;
        pixel_data[0][12] = 0;
        pixel_data[0][13] = 0;
        pixel_data[0][14] = 0;
        pixel_data[0][15] = 0;
        pixel_data[0][16] = 0;
        pixel_data[0][17] = 0;
        pixel_data[0][18] = 0;
        pixel_data[0][19] = 0;
        pixel_data[0][20] = 0;
        pixel_data[0][21] = 0;
        pixel_data[0][22] = 0;
        pixel_data[0][23] = 0;
        pixel_data[0][24] = 0; // y=0
        pixel_data[1][0] = 0;
        pixel_data[1][1] = 0;
        pixel_data[1][2] = 0;
        pixel_data[1][3] = 0;
        pixel_data[1][4] = 0;
        pixel_data[1][5] = 0;
        pixel_data[1][6] = 0;
        pixel_data[1][7] = 0;
        pixel_data[1][8] = 0;
        pixel_data[1][9] = 0;
        pixel_data[1][10] = 0;
        pixel_data[1][11] = 0;
        pixel_data[1][12] = 0;
        pixel_data[1][13] = 0;
        pixel_data[1][14] = 0;
        pixel_data[1][15] = 0;
        pixel_data[1][16] = 0;
        pixel_data[1][17] = 0;
        pixel_data[1][18] = 0;
        pixel_data[1][19] = 0;
        pixel_data[1][20] = 0;
        pixel_data[1][21] = 0;
        pixel_data[1][22] = 0;
        pixel_data[1][23] = 0;
        pixel_data[1][24] = 0; // y=1
        pixel_data[2][0] = 0;
        pixel_data[2][1] = 0;
        pixel_data[2][2] = 0;
        pixel_data[2][3] = 0;
        pixel_data[2][4] = 0;
        pixel_data[2][5] = 0;
        pixel_data[2][6] = 0;
        pixel_data[2][7] = 0;
        pixel_data[2][8] = 0;
        pixel_data[2][9] = 0;
        pixel_data[2][10] = 0;
        pixel_data[2][11] = 0;
        pixel_data[2][12] = 0;
        pixel_data[2][13] = 0;
        pixel_data[2][14] = 0;
        pixel_data[2][15] = 0;
        pixel_data[2][16] = 0;
        pixel_data[2][17] = 0;
        pixel_data[2][18] = 0;
        pixel_data[2][19] = 0;
        pixel_data[2][20] = 0;
        pixel_data[2][21] = 0;
        pixel_data[2][22] = 0;
        pixel_data[2][23] = 0;
        pixel_data[2][24] = 0; // y=2
        pixel_data[3][0] = 0;
        pixel_data[3][1] = 0;
        pixel_data[3][2] = 0;
        pixel_data[3][3] = 0;
        pixel_data[3][4] = 0;
        pixel_data[3][5] = 0;
        pixel_data[3][6] = 0;
        pixel_data[3][7] = 0;
        pixel_data[3][8] = 0;
        pixel_data[3][9] = 0;
        pixel_data[3][10] = 0;
        pixel_data[3][11] = 0;
        pixel_data[3][12] = 0;
        pixel_data[3][13] = 0;
        pixel_data[3][14] = 0;
        pixel_data[3][15] = 0;
        pixel_data[3][16] = 0;
        pixel_data[3][17] = 0;
        pixel_data[3][18] = 0;
        pixel_data[3][19] = 0;
        pixel_data[3][20] = 0;
        pixel_data[3][21] = 0;
        pixel_data[3][22] = 0;
        pixel_data[3][23] = 0;
        pixel_data[3][24] = 0; // y=3
        pixel_data[4][0] = 0;
        pixel_data[4][1] = 0;
        pixel_data[4][2] = 0;
        pixel_data[4][3] = 0;
        pixel_data[4][4] = 0;
        pixel_data[4][5] = 0;
        pixel_data[4][6] = 0;
        pixel_data[4][7] = 0;
        pixel_data[4][8] = 0;
        pixel_data[4][9] = 0;
        pixel_data[4][10] = 0;
        pixel_data[4][11] = 0;
        pixel_data[4][12] = 0;
        pixel_data[4][13] = 0;
        pixel_data[4][14] = 0;
        pixel_data[4][15] = 0;
        pixel_data[4][16] = 0;
        pixel_data[4][17] = 0;
        pixel_data[4][18] = 0;
        pixel_data[4][19] = 0;
        pixel_data[4][20] = 0;
        pixel_data[4][21] = 0;
        pixel_data[4][22] = 0;
        pixel_data[4][23] = 0;
        pixel_data[4][24] = 0; // y=4
        pixel_data[5][0] = 0;
        pixel_data[5][1] = 0;
        pixel_data[5][2] = 0;
        pixel_data[5][3] = 0;
        pixel_data[5][4] = 0;
        pixel_data[5][5] = 0;
        pixel_data[5][6] = 0;
        pixel_data[5][7] = 0;
        pixel_data[5][8] = 0;
        pixel_data[5][9] = 0;
        pixel_data[5][10] = 0;
        pixel_data[5][11] = 0;
        pixel_data[5][12] = 12;
        pixel_data[5][13] = 15;
        pixel_data[5][14] = 14;
        pixel_data[5][15] = 2;
        pixel_data[5][16] = 2;
        pixel_data[5][17] = 2;
        pixel_data[5][18] = 2;
        pixel_data[5][19] = 2;
        pixel_data[5][20] = 15;
        pixel_data[5][21] = 0;
        pixel_data[5][22] = 0;
        pixel_data[5][23] = 0;
        pixel_data[5][24] = 0; // y=5
        pixel_data[6][0] = 0;
        pixel_data[6][1] = 0;
        pixel_data[6][2] = 0;
        pixel_data[6][3] = 0;
        pixel_data[6][4] = 0;
        pixel_data[6][5] = 0;
        pixel_data[6][6] = 0;
        pixel_data[6][7] = 0;
        pixel_data[6][8] = 15;
        pixel_data[6][9] = 14;
        pixel_data[6][10] = 13;
        pixel_data[6][11] = 2;
        pixel_data[6][12] = 0;
        pixel_data[6][13] = 0;
        pixel_data[6][14] = 0;
        pixel_data[6][15] = 0;
        pixel_data[6][16] = 0;
        pixel_data[6][17] = 0;
        pixel_data[6][18] = 0;
        pixel_data[6][19] = 0;
        pixel_data[6][20] = 0;
        pixel_data[6][21] = 15;
        pixel_data[6][22] = 2;
        pixel_data[6][23] = 0;
        pixel_data[6][24] = 0; // y=6
        pixel_data[7][0] = 0;
        pixel_data[7][1] = 0;
        pixel_data[7][2] = 0;
        pixel_data[7][3] = 0;
        pixel_data[7][4] = 14;
        pixel_data[7][5] = 13;
        pixel_data[7][6] = 13;
        pixel_data[7][7] = 15;
        pixel_data[7][8] = 0;
        pixel_data[7][9] = 0;
        pixel_data[7][10] = 0;
        pixel_data[7][11] = 0;
        pixel_data[7][12] = 15;
        pixel_data[7][13] = 15;
        pixel_data[7][14] = 15;
        pixel_data[7][15] = 15;
        pixel_data[7][16] = 15;
        pixel_data[7][17] = 15;
        pixel_data[7][18] = 15;
        pixel_data[7][19] = 15;
        pixel_data[7][20] = 15;
        pixel_data[7][21] = 0;
        pixel_data[7][22] = 0;
        pixel_data[7][23] = 2;
        pixel_data[7][24] = 0; // y=7
        pixel_data[8][0] = 0;
        pixel_data[8][1] = 14;
        pixel_data[8][2] = 2;
        pixel_data[8][3] = 0;
        pixel_data[8][4] = 0;
        pixel_data[8][5] = 0;
        pixel_data[8][6] = 0;
        pixel_data[8][7] = 0;
        pixel_data[8][8] = 15;
        pixel_data[8][9] = 15;
        pixel_data[8][10] = 15;
        pixel_data[8][11] = 15;
        pixel_data[8][12] = 15;
        pixel_data[8][13] = 15;
        pixel_data[8][14] = 15;
        pixel_data[8][15] = 15;
        pixel_data[8][16] = 15;
        pixel_data[8][17] = 15;
        pixel_data[8][18] = 15;
        pixel_data[8][19] = 15;
        pixel_data[8][20] = 15;
        pixel_data[8][21] = 15;
        pixel_data[8][22] = 15;
        pixel_data[8][23] = 0;
        pixel_data[8][24] = 3; // y=8
        pixel_data[9][0] = 14;
        pixel_data[9][1] = 0;
        pixel_data[9][2] = 0;
        pixel_data[9][3] = 15;
        pixel_data[9][4] = 15;
        pixel_data[9][5] = 15;
        pixel_data[9][6] = 15;
        pixel_data[9][7] = 15;
        pixel_data[9][8] = 15;
        pixel_data[9][9] = 15;
        pixel_data[9][10] = 15;
        pixel_data[9][11] = 15;
        pixel_data[9][12] = 15;
        pixel_data[9][13] = 15;
        pixel_data[9][14] = 15;
        pixel_data[9][15] = 15;
        pixel_data[9][16] = 15;
        pixel_data[9][17] = 15;
        pixel_data[9][18] = 15;
        pixel_data[9][19] = 15;
        pixel_data[9][20] = 15;
        pixel_data[9][21] = 15;
        pixel_data[9][22] = 15;
        pixel_data[9][23] = 15;
        pixel_data[9][24] = 0; // y=9
        pixel_data[10][0] = 0;
        pixel_data[10][1] = 15;
        pixel_data[10][2] = 15;
        pixel_data[10][3] = 15;
        pixel_data[10][4] = 15;
        pixel_data[10][5] = 15;
        pixel_data[10][6] = 15;
        pixel_data[10][7] = 15;
        pixel_data[10][8] = 15;
        pixel_data[10][9] = 15;
        pixel_data[10][10] = 15;
        pixel_data[10][11] = 15;
        pixel_data[10][12] = 15;
        pixel_data[10][13] = 15;
        pixel_data[10][14] = 15;
        pixel_data[10][15] = 15;
        pixel_data[10][16] = 15;
        pixel_data[10][17] = 15;
        pixel_data[10][18] = 15;
        pixel_data[10][19] = 15;
        pixel_data[10][20] = 15;
        pixel_data[10][21] = 15;
        pixel_data[10][22] = 15;
        pixel_data[10][23] = 15;
        pixel_data[10][24] = 15; // y=10
        pixel_data[11][0] = 15;
        pixel_data[11][1] = 15;
        pixel_data[11][2] = 15;
        pixel_data[11][3] = 15;
        pixel_data[11][4] = 15;
        pixel_data[11][5] = 15;
        pixel_data[11][6] = 15;
        pixel_data[11][7] = 15;
        pixel_data[11][8] = 15;
        pixel_data[11][9] = 15;
        pixel_data[11][10] = 15;
        pixel_data[11][11] = 15;
        pixel_data[11][12] = 15;
        pixel_data[11][13] = 15;
        pixel_data[11][14] = 15;
        pixel_data[11][15] = 15;
        pixel_data[11][16] = 15;
        pixel_data[11][17] = 15;
        pixel_data[11][18] = 15;
        pixel_data[11][19] = 15;
        pixel_data[11][20] = 15;
        pixel_data[11][21] = 15;
        pixel_data[11][22] = 15;
        pixel_data[11][23] = 15;
        pixel_data[11][24] = 15; // y=11
        pixel_data[12][0] = 15;
        pixel_data[12][1] = 15;
        pixel_data[12][2] = 15;
        pixel_data[12][3] = 15;
        pixel_data[12][4] = 15;
        pixel_data[12][5] = 15;
        pixel_data[12][6] = 15;
        pixel_data[12][7] = 15;
        pixel_data[12][8] = 15;
        pixel_data[12][9] = 15;
        pixel_data[12][10] = 15;
        pixel_data[12][11] = 15;
        pixel_data[12][12] = 15;
        pixel_data[12][13] = 15;
        pixel_data[12][14] = 15;
        pixel_data[12][15] = 15;
        pixel_data[12][16] = 15;
        pixel_data[12][17] = 15;
        pixel_data[12][18] = 15;
        pixel_data[12][19] = 15;
        pixel_data[12][20] = 15;
        pixel_data[12][21] = 15;
        pixel_data[12][22] = 15;
        pixel_data[12][23] = 15;
        pixel_data[12][24] = 15; // y=12
        pixel_data[13][0] = 15;
        pixel_data[13][1] = 15;
        pixel_data[13][2] = 15;
        pixel_data[13][3] = 15;
        pixel_data[13][4] = 15;
        pixel_data[13][5] = 15;
        pixel_data[13][6] = 15;
        pixel_data[13][7] = 15;
        pixel_data[13][8] = 15;
        pixel_data[13][9] = 15;
        pixel_data[13][10] = 15;
        pixel_data[13][11] = 15;
        pixel_data[13][12] = 15;
        pixel_data[13][13] = 15;
        pixel_data[13][14] = 15;
        pixel_data[13][15] = 15;
        pixel_data[13][16] = 15;
        pixel_data[13][17] = 15;
        pixel_data[13][18] = 15;
        pixel_data[13][19] = 15;
        pixel_data[13][20] = 15;
        pixel_data[13][21] = 15;
        pixel_data[13][22] = 15;
        pixel_data[13][23] = 15;
        pixel_data[13][24] = 15; // y=13
        pixel_data[14][0] = 0;
        pixel_data[14][1] = 15;
        pixel_data[14][2] = 15;
        pixel_data[14][3] = 15;
        pixel_data[14][4] = 15;
        pixel_data[14][5] = 15;
        pixel_data[14][6] = 15;
        pixel_data[14][7] = 15;
        pixel_data[14][8] = 15;
        pixel_data[14][9] = 15;
        pixel_data[14][10] = 15;
        pixel_data[14][11] = 15;
        pixel_data[14][12] = 15;
        pixel_data[14][13] = 1;
        pixel_data[14][14] = 1;
        pixel_data[14][15] = 15;
        pixel_data[14][16] = 15;
        pixel_data[14][17] = 15;
        pixel_data[14][18] = 15;
        pixel_data[14][19] = 15;
        pixel_data[14][20] = 15;
        pixel_data[14][21] = 15;
        pixel_data[14][22] = 15;
        pixel_data[14][23] = 15;
        pixel_data[14][24] = 15; // y=14
        pixel_data[15][0] = 2;
        pixel_data[15][1] = 0;
        pixel_data[15][2] = 0;
        pixel_data[15][3] = 0;
        pixel_data[15][4] = 0;
        pixel_data[15][5] = 0;
        pixel_data[15][6] = 0;
        pixel_data[15][7] = 13;
        pixel_data[15][8] = 15;
        pixel_data[15][9] = 15;
        pixel_data[15][10] = 15;
        pixel_data[15][11] = 15;
        pixel_data[15][12] = 15;
        pixel_data[15][13] = 15;
        pixel_data[15][14] = 15;
        pixel_data[15][15] = 15;
        pixel_data[15][16] = 15;
        pixel_data[15][17] = 15;
        pixel_data[15][18] = 15;
        pixel_data[15][19] = 15;
        pixel_data[15][20] = 15;
        pixel_data[15][21] = 15;
        pixel_data[15][22] = 15;
        pixel_data[15][23] = 13;
        pixel_data[15][24] = 0; // y=15
        pixel_data[16][0] = 0;
        pixel_data[16][1] = 15;
        pixel_data[16][2] = 13;
        pixel_data[16][3] = 3;
        pixel_data[16][4] = 15;
        pixel_data[16][5] = 13;
        pixel_data[16][6] = 15;
        pixel_data[16][7] = 0;
        pixel_data[16][8] = 0;
        pixel_data[16][9] = 0;
        pixel_data[16][10] = 0;
        pixel_data[16][11] = 0;
        pixel_data[16][12] = 0;
        pixel_data[16][13] = 0;
        pixel_data[16][14] = 0;
        pixel_data[16][15] = 4;
        pixel_data[16][16] = 15;
        pixel_data[16][17] = 15;
        pixel_data[16][18] = 15;
        pixel_data[16][19] = 15;
        pixel_data[16][20] = 15;
        pixel_data[16][21] = 0;
        pixel_data[16][22] = 0;
        pixel_data[16][23] = 0;
        pixel_data[16][24] = 14; // y=16
        pixel_data[17][0] = 0;
        pixel_data[17][1] = 0;
        pixel_data[17][2] = 0;
        pixel_data[17][3] = 0;
        pixel_data[17][4] = 0;
        pixel_data[17][5] = 0;
        pixel_data[17][6] = 0;
        pixel_data[17][7] = 15;
        pixel_data[17][8] = 15;
        pixel_data[17][9] = 2;
        pixel_data[17][10] = 13;
        pixel_data[17][11] = 15;
        pixel_data[17][12] = 15;
        pixel_data[17][13] = 15;
        pixel_data[17][14] = 0;
        pixel_data[17][15] = 0;
        pixel_data[17][16] = 0;
        pixel_data[17][17] = 0;
        pixel_data[17][18] = 0;
        pixel_data[17][19] = 0;
        pixel_data[17][20] = 0;
        pixel_data[17][21] = 2;
        pixel_data[17][22] = 4;
        pixel_data[17][23] = 15;
        pixel_data[17][24] = 0; // y=17
        pixel_data[18][0] = 0;
        pixel_data[18][1] = 0;
        pixel_data[18][2] = 0;
        pixel_data[18][3] = 0;
        pixel_data[18][4] = 0;
        pixel_data[18][5] = 0;
        pixel_data[18][6] = 0;
        pixel_data[18][7] = 0;
        pixel_data[18][8] = 0;
        pixel_data[18][9] = 0;
        pixel_data[18][10] = 0;
        pixel_data[18][11] = 0;
        pixel_data[18][12] = 0;
        pixel_data[18][13] = 0;
        pixel_data[18][14] = 0;
        pixel_data[18][15] = 15;
        pixel_data[18][16] = 3;
        pixel_data[18][17] = 13;
        pixel_data[18][18] = 13;
        pixel_data[18][19] = 13;
        pixel_data[18][20] = 15;
        pixel_data[18][21] = 0;
        pixel_data[18][22] = 0;
        pixel_data[18][23] = 0;
        pixel_data[18][24] = 0; // y=18
        pixel_data[19][0] = 0;
        pixel_data[19][1] = 0;
        pixel_data[19][2] = 0;
        pixel_data[19][3] = 0;
        pixel_data[19][4] = 0;
        pixel_data[19][5] = 0;
        pixel_data[19][6] = 0;
        pixel_data[19][7] = 0;
        pixel_data[19][8] = 0;
        pixel_data[19][9] = 0;
        pixel_data[19][10] = 0;
        pixel_data[19][11] = 0;
        pixel_data[19][12] = 0;
        pixel_data[19][13] = 0;
        pixel_data[19][14] = 0;
        pixel_data[19][15] = 0;
        pixel_data[19][16] = 0;
        pixel_data[19][17] = 0;
        pixel_data[19][18] = 0;
        pixel_data[19][19] = 0;
        pixel_data[19][20] = 0;
        pixel_data[19][21] = 0;
        pixel_data[19][22] = 0;
        pixel_data[19][23] = 0;
        pixel_data[19][24] = 0; // y=19
        pixel_data[20][0] = 0;
        pixel_data[20][1] = 0;
        pixel_data[20][2] = 0;
        pixel_data[20][3] = 0;
        pixel_data[20][4] = 0;
        pixel_data[20][5] = 0;
        pixel_data[20][6] = 0;
        pixel_data[20][7] = 0;
        pixel_data[20][8] = 0;
        pixel_data[20][9] = 0;
        pixel_data[20][10] = 0;
        pixel_data[20][11] = 0;
        pixel_data[20][12] = 0;
        pixel_data[20][13] = 0;
        pixel_data[20][14] = 0;
        pixel_data[20][15] = 0;
        pixel_data[20][16] = 0;
        pixel_data[20][17] = 0;
        pixel_data[20][18] = 0;
        pixel_data[20][19] = 0;
        pixel_data[20][20] = 0;
        pixel_data[20][21] = 0;
        pixel_data[20][22] = 0;
        pixel_data[20][23] = 0;
        pixel_data[20][24] = 0; // y=20
        pixel_data[21][0] = 0;
        pixel_data[21][1] = 0;
        pixel_data[21][2] = 0;
        pixel_data[21][3] = 0;
        pixel_data[21][4] = 0;
        pixel_data[21][5] = 0;
        pixel_data[21][6] = 0;
        pixel_data[21][7] = 0;
        pixel_data[21][8] = 0;
        pixel_data[21][9] = 0;
        pixel_data[21][10] = 0;
        pixel_data[21][11] = 0;
        pixel_data[21][12] = 0;
        pixel_data[21][13] = 0;
        pixel_data[21][14] = 0;
        pixel_data[21][15] = 0;
        pixel_data[21][16] = 0;
        pixel_data[21][17] = 0;
        pixel_data[21][18] = 0;
        pixel_data[21][19] = 0;
        pixel_data[21][20] = 0;
        pixel_data[21][21] = 0;
        pixel_data[21][22] = 0;
        pixel_data[21][23] = 0;
        pixel_data[21][24] = 0; // y=21
        pixel_data[22][0] = 0;
        pixel_data[22][1] = 0;
        pixel_data[22][2] = 0;
        pixel_data[22][3] = 0;
        pixel_data[22][4] = 0;
        pixel_data[22][5] = 0;
        pixel_data[22][6] = 0;
        pixel_data[22][7] = 0;
        pixel_data[22][8] = 0;
        pixel_data[22][9] = 0;
        pixel_data[22][10] = 0;
        pixel_data[22][11] = 0;
        pixel_data[22][12] = 0;
        pixel_data[22][13] = 0;
        pixel_data[22][14] = 0;
        pixel_data[22][15] = 0;
        pixel_data[22][16] = 0;
        pixel_data[22][17] = 0;
        pixel_data[22][18] = 0;
        pixel_data[22][19] = 0;
        pixel_data[22][20] = 0;
        pixel_data[22][21] = 0;
        pixel_data[22][22] = 0;
        pixel_data[22][23] = 0;
        pixel_data[22][24] = 0; // y=22
        pixel_data[23][0] = 0;
        pixel_data[23][1] = 0;
        pixel_data[23][2] = 0;
        pixel_data[23][3] = 0;
        pixel_data[23][4] = 0;
        pixel_data[23][5] = 0;
        pixel_data[23][6] = 0;
        pixel_data[23][7] = 0;
        pixel_data[23][8] = 0;
        pixel_data[23][9] = 0;
        pixel_data[23][10] = 0;
        pixel_data[23][11] = 0;
        pixel_data[23][12] = 0;
        pixel_data[23][13] = 0;
        pixel_data[23][14] = 0;
        pixel_data[23][15] = 0;
        pixel_data[23][16] = 0;
        pixel_data[23][17] = 0;
        pixel_data[23][18] = 0;
        pixel_data[23][19] = 0;
        pixel_data[23][20] = 0;
        pixel_data[23][21] = 0;
        pixel_data[23][22] = 0;
        pixel_data[23][23] = 0;
        pixel_data[23][24] = 0; // y=23
        pixel_data[24][0] = 0;
        pixel_data[24][1] = 0;
        pixel_data[24][2] = 0;
        pixel_data[24][3] = 0;
        pixel_data[24][4] = 0;
        pixel_data[24][5] = 0;
        pixel_data[24][6] = 0;
        pixel_data[24][7] = 0;
        pixel_data[24][8] = 0;
        pixel_data[24][9] = 0;
        pixel_data[24][10] = 0;
        pixel_data[24][11] = 0;
        pixel_data[24][12] = 0;
        pixel_data[24][13] = 0;
        pixel_data[24][14] = 0;
        pixel_data[24][15] = 0;
        pixel_data[24][16] = 0;
        pixel_data[24][17] = 0;
        pixel_data[24][18] = 0;
        pixel_data[24][19] = 0;
        pixel_data[24][20] = 0;
        pixel_data[24][21] = 0;
        pixel_data[24][22] = 0;
        pixel_data[24][23] = 0;
        pixel_data[24][24] = 0; // y=24
    end
endmodule
