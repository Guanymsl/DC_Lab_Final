module player1_squat_lut(output reg [3:0] pixel_data [0:199][0:199]);
    initial begin
        pixel_data[0][0] = 0;
        pixel_data[0][1] = 0;
        pixel_data[0][2] = 0;
        pixel_data[0][3] = 0;
        pixel_data[0][4] = 0;
        pixel_data[0][5] = 0;
        pixel_data[0][6] = 0;
        pixel_data[0][7] = 0;
        pixel_data[0][8] = 0;
        pixel_data[0][9] = 0;
        pixel_data[0][10] = 0;
        pixel_data[0][11] = 0;
        pixel_data[0][12] = 0;
        pixel_data[0][13] = 0;
        pixel_data[0][14] = 0;
        pixel_data[0][15] = 0;
        pixel_data[0][16] = 0;
        pixel_data[0][17] = 0;
        pixel_data[0][18] = 0;
        pixel_data[0][19] = 0;
        pixel_data[0][20] = 0;
        pixel_data[0][21] = 0;
        pixel_data[0][22] = 0;
        pixel_data[0][23] = 0;
        pixel_data[0][24] = 0;
        pixel_data[0][25] = 0;
        pixel_data[0][26] = 0;
        pixel_data[0][27] = 0;
        pixel_data[0][28] = 0;
        pixel_data[0][29] = 0;
        pixel_data[0][30] = 0;
        pixel_data[0][31] = 0;
        pixel_data[0][32] = 0;
        pixel_data[0][33] = 0;
        pixel_data[0][34] = 0;
        pixel_data[0][35] = 0;
        pixel_data[0][36] = 0;
        pixel_data[0][37] = 0;
        pixel_data[0][38] = 0;
        pixel_data[0][39] = 0;
        pixel_data[0][40] = 0;
        pixel_data[0][41] = 0;
        pixel_data[0][42] = 0;
        pixel_data[0][43] = 0;
        pixel_data[0][44] = 0;
        pixel_data[0][45] = 0;
        pixel_data[0][46] = 0;
        pixel_data[0][47] = 0;
        pixel_data[0][48] = 0;
        pixel_data[0][49] = 0;
        pixel_data[0][50] = 0;
        pixel_data[0][51] = 0;
        pixel_data[0][52] = 0;
        pixel_data[0][53] = 0;
        pixel_data[0][54] = 0;
        pixel_data[0][55] = 0;
        pixel_data[0][56] = 0;
        pixel_data[0][57] = 0;
        pixel_data[0][58] = 0;
        pixel_data[0][59] = 0;
        pixel_data[0][60] = 0;
        pixel_data[0][61] = 0;
        pixel_data[0][62] = 0;
        pixel_data[0][63] = 0;
        pixel_data[0][64] = 0;
        pixel_data[0][65] = 0;
        pixel_data[0][66] = 0;
        pixel_data[0][67] = 0;
        pixel_data[0][68] = 0;
        pixel_data[0][69] = 0;
        pixel_data[0][70] = 0;
        pixel_data[0][71] = 0;
        pixel_data[0][72] = 0;
        pixel_data[0][73] = 0;
        pixel_data[0][74] = 0;
        pixel_data[0][75] = 0;
        pixel_data[0][76] = 0;
        pixel_data[0][77] = 0;
        pixel_data[0][78] = 0;
        pixel_data[0][79] = 0;
        pixel_data[0][80] = 0;
        pixel_data[0][81] = 0;
        pixel_data[0][82] = 0;
        pixel_data[0][83] = 0;
        pixel_data[0][84] = 0;
        pixel_data[0][85] = 0;
        pixel_data[0][86] = 0;
        pixel_data[0][87] = 0;
        pixel_data[0][88] = 0;
        pixel_data[0][89] = 0;
        pixel_data[0][90] = 0;
        pixel_data[0][91] = 0;
        pixel_data[0][92] = 0;
        pixel_data[0][93] = 0;
        pixel_data[0][94] = 0;
        pixel_data[0][95] = 0;
        pixel_data[0][96] = 0;
        pixel_data[0][97] = 0;
        pixel_data[0][98] = 0;
        pixel_data[0][99] = 0;
        pixel_data[0][100] = 0;
        pixel_data[0][101] = 0;
        pixel_data[0][102] = 0;
        pixel_data[0][103] = 0;
        pixel_data[0][104] = 0;
        pixel_data[0][105] = 0;
        pixel_data[0][106] = 0;
        pixel_data[0][107] = 0;
        pixel_data[0][108] = 0;
        pixel_data[0][109] = 0;
        pixel_data[0][110] = 0;
        pixel_data[0][111] = 0;
        pixel_data[0][112] = 0;
        pixel_data[0][113] = 0;
        pixel_data[0][114] = 0;
        pixel_data[0][115] = 0;
        pixel_data[0][116] = 0;
        pixel_data[0][117] = 0;
        pixel_data[0][118] = 0;
        pixel_data[0][119] = 0;
        pixel_data[0][120] = 0;
        pixel_data[0][121] = 0;
        pixel_data[0][122] = 0;
        pixel_data[0][123] = 0;
        pixel_data[0][124] = 0;
        pixel_data[0][125] = 0;
        pixel_data[0][126] = 0;
        pixel_data[0][127] = 0;
        pixel_data[0][128] = 0;
        pixel_data[0][129] = 0;
        pixel_data[0][130] = 0;
        pixel_data[0][131] = 0;
        pixel_data[0][132] = 0;
        pixel_data[0][133] = 0;
        pixel_data[0][134] = 0;
        pixel_data[0][135] = 0;
        pixel_data[0][136] = 0;
        pixel_data[0][137] = 0;
        pixel_data[0][138] = 0;
        pixel_data[0][139] = 0;
        pixel_data[0][140] = 0;
        pixel_data[0][141] = 0;
        pixel_data[0][142] = 0;
        pixel_data[0][143] = 0;
        pixel_data[0][144] = 0;
        pixel_data[0][145] = 0;
        pixel_data[0][146] = 0;
        pixel_data[0][147] = 0;
        pixel_data[0][148] = 0;
        pixel_data[0][149] = 0;
        pixel_data[0][150] = 0;
        pixel_data[0][151] = 0;
        pixel_data[0][152] = 0;
        pixel_data[0][153] = 0;
        pixel_data[0][154] = 0;
        pixel_data[0][155] = 0;
        pixel_data[0][156] = 0;
        pixel_data[0][157] = 0;
        pixel_data[0][158] = 0;
        pixel_data[0][159] = 0;
        pixel_data[0][160] = 0;
        pixel_data[0][161] = 0;
        pixel_data[0][162] = 0;
        pixel_data[0][163] = 0;
        pixel_data[0][164] = 0;
        pixel_data[0][165] = 0;
        pixel_data[0][166] = 0;
        pixel_data[0][167] = 0;
        pixel_data[0][168] = 0;
        pixel_data[0][169] = 0;
        pixel_data[0][170] = 0;
        pixel_data[0][171] = 0;
        pixel_data[0][172] = 0;
        pixel_data[0][173] = 0;
        pixel_data[0][174] = 0;
        pixel_data[0][175] = 0;
        pixel_data[0][176] = 0;
        pixel_data[0][177] = 0;
        pixel_data[0][178] = 0;
        pixel_data[0][179] = 0;
        pixel_data[0][180] = 0;
        pixel_data[0][181] = 0;
        pixel_data[0][182] = 0;
        pixel_data[0][183] = 0;
        pixel_data[0][184] = 0;
        pixel_data[0][185] = 0;
        pixel_data[0][186] = 0;
        pixel_data[0][187] = 0;
        pixel_data[0][188] = 0;
        pixel_data[0][189] = 0;
        pixel_data[0][190] = 0;
        pixel_data[0][191] = 0;
        pixel_data[0][192] = 0;
        pixel_data[0][193] = 0;
        pixel_data[0][194] = 0;
        pixel_data[0][195] = 0;
        pixel_data[0][196] = 0;
        pixel_data[0][197] = 0;
        pixel_data[0][198] = 0;
        pixel_data[0][199] = 0; // y=0
        pixel_data[1][0] = 0;
        pixel_data[1][1] = 0;
        pixel_data[1][2] = 0;
        pixel_data[1][3] = 0;
        pixel_data[1][4] = 0;
        pixel_data[1][5] = 0;
        pixel_data[1][6] = 0;
        pixel_data[1][7] = 0;
        pixel_data[1][8] = 0;
        pixel_data[1][9] = 0;
        pixel_data[1][10] = 0;
        pixel_data[1][11] = 0;
        pixel_data[1][12] = 0;
        pixel_data[1][13] = 0;
        pixel_data[1][14] = 0;
        pixel_data[1][15] = 0;
        pixel_data[1][16] = 0;
        pixel_data[1][17] = 0;
        pixel_data[1][18] = 0;
        pixel_data[1][19] = 0;
        pixel_data[1][20] = 0;
        pixel_data[1][21] = 0;
        pixel_data[1][22] = 0;
        pixel_data[1][23] = 0;
        pixel_data[1][24] = 0;
        pixel_data[1][25] = 0;
        pixel_data[1][26] = 0;
        pixel_data[1][27] = 0;
        pixel_data[1][28] = 0;
        pixel_data[1][29] = 0;
        pixel_data[1][30] = 0;
        pixel_data[1][31] = 0;
        pixel_data[1][32] = 0;
        pixel_data[1][33] = 0;
        pixel_data[1][34] = 0;
        pixel_data[1][35] = 0;
        pixel_data[1][36] = 0;
        pixel_data[1][37] = 0;
        pixel_data[1][38] = 0;
        pixel_data[1][39] = 0;
        pixel_data[1][40] = 0;
        pixel_data[1][41] = 0;
        pixel_data[1][42] = 0;
        pixel_data[1][43] = 0;
        pixel_data[1][44] = 0;
        pixel_data[1][45] = 0;
        pixel_data[1][46] = 0;
        pixel_data[1][47] = 0;
        pixel_data[1][48] = 0;
        pixel_data[1][49] = 0;
        pixel_data[1][50] = 0;
        pixel_data[1][51] = 0;
        pixel_data[1][52] = 0;
        pixel_data[1][53] = 0;
        pixel_data[1][54] = 0;
        pixel_data[1][55] = 0;
        pixel_data[1][56] = 0;
        pixel_data[1][57] = 0;
        pixel_data[1][58] = 0;
        pixel_data[1][59] = 0;
        pixel_data[1][60] = 0;
        pixel_data[1][61] = 0;
        pixel_data[1][62] = 0;
        pixel_data[1][63] = 0;
        pixel_data[1][64] = 0;
        pixel_data[1][65] = 0;
        pixel_data[1][66] = 0;
        pixel_data[1][67] = 0;
        pixel_data[1][68] = 0;
        pixel_data[1][69] = 0;
        pixel_data[1][70] = 0;
        pixel_data[1][71] = 0;
        pixel_data[1][72] = 0;
        pixel_data[1][73] = 0;
        pixel_data[1][74] = 0;
        pixel_data[1][75] = 0;
        pixel_data[1][76] = 0;
        pixel_data[1][77] = 0;
        pixel_data[1][78] = 0;
        pixel_data[1][79] = 0;
        pixel_data[1][80] = 0;
        pixel_data[1][81] = 0;
        pixel_data[1][82] = 0;
        pixel_data[1][83] = 0;
        pixel_data[1][84] = 0;
        pixel_data[1][85] = 0;
        pixel_data[1][86] = 0;
        pixel_data[1][87] = 0;
        pixel_data[1][88] = 0;
        pixel_data[1][89] = 0;
        pixel_data[1][90] = 0;
        pixel_data[1][91] = 0;
        pixel_data[1][92] = 0;
        pixel_data[1][93] = 0;
        pixel_data[1][94] = 0;
        pixel_data[1][95] = 0;
        pixel_data[1][96] = 0;
        pixel_data[1][97] = 0;
        pixel_data[1][98] = 0;
        pixel_data[1][99] = 0;
        pixel_data[1][100] = 0;
        pixel_data[1][101] = 0;
        pixel_data[1][102] = 0;
        pixel_data[1][103] = 0;
        pixel_data[1][104] = 0;
        pixel_data[1][105] = 0;
        pixel_data[1][106] = 0;
        pixel_data[1][107] = 0;
        pixel_data[1][108] = 0;
        pixel_data[1][109] = 0;
        pixel_data[1][110] = 0;
        pixel_data[1][111] = 0;
        pixel_data[1][112] = 0;
        pixel_data[1][113] = 0;
        pixel_data[1][114] = 0;
        pixel_data[1][115] = 0;
        pixel_data[1][116] = 0;
        pixel_data[1][117] = 0;
        pixel_data[1][118] = 0;
        pixel_data[1][119] = 0;
        pixel_data[1][120] = 0;
        pixel_data[1][121] = 0;
        pixel_data[1][122] = 0;
        pixel_data[1][123] = 0;
        pixel_data[1][124] = 0;
        pixel_data[1][125] = 0;
        pixel_data[1][126] = 0;
        pixel_data[1][127] = 0;
        pixel_data[1][128] = 0;
        pixel_data[1][129] = 0;
        pixel_data[1][130] = 0;
        pixel_data[1][131] = 0;
        pixel_data[1][132] = 0;
        pixel_data[1][133] = 0;
        pixel_data[1][134] = 0;
        pixel_data[1][135] = 0;
        pixel_data[1][136] = 0;
        pixel_data[1][137] = 0;
        pixel_data[1][138] = 0;
        pixel_data[1][139] = 0;
        pixel_data[1][140] = 0;
        pixel_data[1][141] = 0;
        pixel_data[1][142] = 0;
        pixel_data[1][143] = 0;
        pixel_data[1][144] = 0;
        pixel_data[1][145] = 0;
        pixel_data[1][146] = 0;
        pixel_data[1][147] = 0;
        pixel_data[1][148] = 0;
        pixel_data[1][149] = 0;
        pixel_data[1][150] = 0;
        pixel_data[1][151] = 0;
        pixel_data[1][152] = 0;
        pixel_data[1][153] = 0;
        pixel_data[1][154] = 0;
        pixel_data[1][155] = 0;
        pixel_data[1][156] = 0;
        pixel_data[1][157] = 0;
        pixel_data[1][158] = 0;
        pixel_data[1][159] = 0;
        pixel_data[1][160] = 0;
        pixel_data[1][161] = 0;
        pixel_data[1][162] = 0;
        pixel_data[1][163] = 0;
        pixel_data[1][164] = 0;
        pixel_data[1][165] = 0;
        pixel_data[1][166] = 0;
        pixel_data[1][167] = 0;
        pixel_data[1][168] = 0;
        pixel_data[1][169] = 0;
        pixel_data[1][170] = 0;
        pixel_data[1][171] = 0;
        pixel_data[1][172] = 0;
        pixel_data[1][173] = 0;
        pixel_data[1][174] = 0;
        pixel_data[1][175] = 0;
        pixel_data[1][176] = 0;
        pixel_data[1][177] = 0;
        pixel_data[1][178] = 0;
        pixel_data[1][179] = 0;
        pixel_data[1][180] = 0;
        pixel_data[1][181] = 0;
        pixel_data[1][182] = 0;
        pixel_data[1][183] = 0;
        pixel_data[1][184] = 0;
        pixel_data[1][185] = 0;
        pixel_data[1][186] = 0;
        pixel_data[1][187] = 0;
        pixel_data[1][188] = 0;
        pixel_data[1][189] = 0;
        pixel_data[1][190] = 0;
        pixel_data[1][191] = 0;
        pixel_data[1][192] = 0;
        pixel_data[1][193] = 0;
        pixel_data[1][194] = 0;
        pixel_data[1][195] = 0;
        pixel_data[1][196] = 0;
        pixel_data[1][197] = 0;
        pixel_data[1][198] = 0;
        pixel_data[1][199] = 0; // y=1
        pixel_data[2][0] = 0;
        pixel_data[2][1] = 0;
        pixel_data[2][2] = 0;
        pixel_data[2][3] = 0;
        pixel_data[2][4] = 0;
        pixel_data[2][5] = 0;
        pixel_data[2][6] = 0;
        pixel_data[2][7] = 0;
        pixel_data[2][8] = 0;
        pixel_data[2][9] = 0;
        pixel_data[2][10] = 0;
        pixel_data[2][11] = 0;
        pixel_data[2][12] = 0;
        pixel_data[2][13] = 0;
        pixel_data[2][14] = 0;
        pixel_data[2][15] = 0;
        pixel_data[2][16] = 0;
        pixel_data[2][17] = 0;
        pixel_data[2][18] = 0;
        pixel_data[2][19] = 0;
        pixel_data[2][20] = 0;
        pixel_data[2][21] = 0;
        pixel_data[2][22] = 0;
        pixel_data[2][23] = 0;
        pixel_data[2][24] = 0;
        pixel_data[2][25] = 0;
        pixel_data[2][26] = 0;
        pixel_data[2][27] = 0;
        pixel_data[2][28] = 0;
        pixel_data[2][29] = 0;
        pixel_data[2][30] = 0;
        pixel_data[2][31] = 0;
        pixel_data[2][32] = 0;
        pixel_data[2][33] = 0;
        pixel_data[2][34] = 0;
        pixel_data[2][35] = 0;
        pixel_data[2][36] = 0;
        pixel_data[2][37] = 0;
        pixel_data[2][38] = 0;
        pixel_data[2][39] = 0;
        pixel_data[2][40] = 0;
        pixel_data[2][41] = 0;
        pixel_data[2][42] = 0;
        pixel_data[2][43] = 0;
        pixel_data[2][44] = 0;
        pixel_data[2][45] = 0;
        pixel_data[2][46] = 0;
        pixel_data[2][47] = 0;
        pixel_data[2][48] = 0;
        pixel_data[2][49] = 0;
        pixel_data[2][50] = 0;
        pixel_data[2][51] = 0;
        pixel_data[2][52] = 0;
        pixel_data[2][53] = 0;
        pixel_data[2][54] = 0;
        pixel_data[2][55] = 0;
        pixel_data[2][56] = 0;
        pixel_data[2][57] = 0;
        pixel_data[2][58] = 0;
        pixel_data[2][59] = 0;
        pixel_data[2][60] = 0;
        pixel_data[2][61] = 0;
        pixel_data[2][62] = 0;
        pixel_data[2][63] = 0;
        pixel_data[2][64] = 0;
        pixel_data[2][65] = 0;
        pixel_data[2][66] = 0;
        pixel_data[2][67] = 0;
        pixel_data[2][68] = 0;
        pixel_data[2][69] = 0;
        pixel_data[2][70] = 0;
        pixel_data[2][71] = 0;
        pixel_data[2][72] = 0;
        pixel_data[2][73] = 0;
        pixel_data[2][74] = 0;
        pixel_data[2][75] = 0;
        pixel_data[2][76] = 0;
        pixel_data[2][77] = 0;
        pixel_data[2][78] = 0;
        pixel_data[2][79] = 0;
        pixel_data[2][80] = 0;
        pixel_data[2][81] = 0;
        pixel_data[2][82] = 0;
        pixel_data[2][83] = 0;
        pixel_data[2][84] = 0;
        pixel_data[2][85] = 0;
        pixel_data[2][86] = 0;
        pixel_data[2][87] = 0;
        pixel_data[2][88] = 0;
        pixel_data[2][89] = 0;
        pixel_data[2][90] = 0;
        pixel_data[2][91] = 0;
        pixel_data[2][92] = 0;
        pixel_data[2][93] = 0;
        pixel_data[2][94] = 0;
        pixel_data[2][95] = 0;
        pixel_data[2][96] = 0;
        pixel_data[2][97] = 0;
        pixel_data[2][98] = 0;
        pixel_data[2][99] = 0;
        pixel_data[2][100] = 0;
        pixel_data[2][101] = 0;
        pixel_data[2][102] = 0;
        pixel_data[2][103] = 0;
        pixel_data[2][104] = 0;
        pixel_data[2][105] = 0;
        pixel_data[2][106] = 0;
        pixel_data[2][107] = 0;
        pixel_data[2][108] = 0;
        pixel_data[2][109] = 0;
        pixel_data[2][110] = 0;
        pixel_data[2][111] = 0;
        pixel_data[2][112] = 0;
        pixel_data[2][113] = 0;
        pixel_data[2][114] = 0;
        pixel_data[2][115] = 0;
        pixel_data[2][116] = 0;
        pixel_data[2][117] = 0;
        pixel_data[2][118] = 0;
        pixel_data[2][119] = 0;
        pixel_data[2][120] = 0;
        pixel_data[2][121] = 0;
        pixel_data[2][122] = 0;
        pixel_data[2][123] = 0;
        pixel_data[2][124] = 0;
        pixel_data[2][125] = 0;
        pixel_data[2][126] = 0;
        pixel_data[2][127] = 0;
        pixel_data[2][128] = 0;
        pixel_data[2][129] = 0;
        pixel_data[2][130] = 0;
        pixel_data[2][131] = 0;
        pixel_data[2][132] = 0;
        pixel_data[2][133] = 0;
        pixel_data[2][134] = 0;
        pixel_data[2][135] = 0;
        pixel_data[2][136] = 0;
        pixel_data[2][137] = 0;
        pixel_data[2][138] = 0;
        pixel_data[2][139] = 0;
        pixel_data[2][140] = 0;
        pixel_data[2][141] = 0;
        pixel_data[2][142] = 0;
        pixel_data[2][143] = 0;
        pixel_data[2][144] = 0;
        pixel_data[2][145] = 0;
        pixel_data[2][146] = 0;
        pixel_data[2][147] = 0;
        pixel_data[2][148] = 0;
        pixel_data[2][149] = 0;
        pixel_data[2][150] = 0;
        pixel_data[2][151] = 0;
        pixel_data[2][152] = 0;
        pixel_data[2][153] = 0;
        pixel_data[2][154] = 0;
        pixel_data[2][155] = 0;
        pixel_data[2][156] = 0;
        pixel_data[2][157] = 0;
        pixel_data[2][158] = 0;
        pixel_data[2][159] = 0;
        pixel_data[2][160] = 0;
        pixel_data[2][161] = 0;
        pixel_data[2][162] = 0;
        pixel_data[2][163] = 0;
        pixel_data[2][164] = 0;
        pixel_data[2][165] = 0;
        pixel_data[2][166] = 0;
        pixel_data[2][167] = 0;
        pixel_data[2][168] = 0;
        pixel_data[2][169] = 0;
        pixel_data[2][170] = 0;
        pixel_data[2][171] = 0;
        pixel_data[2][172] = 0;
        pixel_data[2][173] = 0;
        pixel_data[2][174] = 0;
        pixel_data[2][175] = 0;
        pixel_data[2][176] = 0;
        pixel_data[2][177] = 0;
        pixel_data[2][178] = 0;
        pixel_data[2][179] = 0;
        pixel_data[2][180] = 0;
        pixel_data[2][181] = 0;
        pixel_data[2][182] = 0;
        pixel_data[2][183] = 0;
        pixel_data[2][184] = 0;
        pixel_data[2][185] = 0;
        pixel_data[2][186] = 0;
        pixel_data[2][187] = 0;
        pixel_data[2][188] = 0;
        pixel_data[2][189] = 0;
        pixel_data[2][190] = 0;
        pixel_data[2][191] = 0;
        pixel_data[2][192] = 0;
        pixel_data[2][193] = 0;
        pixel_data[2][194] = 0;
        pixel_data[2][195] = 0;
        pixel_data[2][196] = 0;
        pixel_data[2][197] = 0;
        pixel_data[2][198] = 0;
        pixel_data[2][199] = 0; // y=2
        pixel_data[3][0] = 0;
        pixel_data[3][1] = 0;
        pixel_data[3][2] = 0;
        pixel_data[3][3] = 0;
        pixel_data[3][4] = 0;
        pixel_data[3][5] = 0;
        pixel_data[3][6] = 0;
        pixel_data[3][7] = 0;
        pixel_data[3][8] = 0;
        pixel_data[3][9] = 0;
        pixel_data[3][10] = 0;
        pixel_data[3][11] = 0;
        pixel_data[3][12] = 0;
        pixel_data[3][13] = 0;
        pixel_data[3][14] = 0;
        pixel_data[3][15] = 0;
        pixel_data[3][16] = 0;
        pixel_data[3][17] = 0;
        pixel_data[3][18] = 0;
        pixel_data[3][19] = 0;
        pixel_data[3][20] = 0;
        pixel_data[3][21] = 0;
        pixel_data[3][22] = 0;
        pixel_data[3][23] = 0;
        pixel_data[3][24] = 0;
        pixel_data[3][25] = 0;
        pixel_data[3][26] = 0;
        pixel_data[3][27] = 0;
        pixel_data[3][28] = 0;
        pixel_data[3][29] = 0;
        pixel_data[3][30] = 0;
        pixel_data[3][31] = 0;
        pixel_data[3][32] = 0;
        pixel_data[3][33] = 0;
        pixel_data[3][34] = 0;
        pixel_data[3][35] = 0;
        pixel_data[3][36] = 0;
        pixel_data[3][37] = 0;
        pixel_data[3][38] = 0;
        pixel_data[3][39] = 0;
        pixel_data[3][40] = 0;
        pixel_data[3][41] = 0;
        pixel_data[3][42] = 0;
        pixel_data[3][43] = 0;
        pixel_data[3][44] = 0;
        pixel_data[3][45] = 0;
        pixel_data[3][46] = 0;
        pixel_data[3][47] = 0;
        pixel_data[3][48] = 0;
        pixel_data[3][49] = 0;
        pixel_data[3][50] = 0;
        pixel_data[3][51] = 0;
        pixel_data[3][52] = 0;
        pixel_data[3][53] = 0;
        pixel_data[3][54] = 0;
        pixel_data[3][55] = 0;
        pixel_data[3][56] = 0;
        pixel_data[3][57] = 0;
        pixel_data[3][58] = 0;
        pixel_data[3][59] = 0;
        pixel_data[3][60] = 0;
        pixel_data[3][61] = 0;
        pixel_data[3][62] = 0;
        pixel_data[3][63] = 0;
        pixel_data[3][64] = 0;
        pixel_data[3][65] = 0;
        pixel_data[3][66] = 0;
        pixel_data[3][67] = 0;
        pixel_data[3][68] = 0;
        pixel_data[3][69] = 0;
        pixel_data[3][70] = 0;
        pixel_data[3][71] = 0;
        pixel_data[3][72] = 0;
        pixel_data[3][73] = 0;
        pixel_data[3][74] = 0;
        pixel_data[3][75] = 0;
        pixel_data[3][76] = 0;
        pixel_data[3][77] = 0;
        pixel_data[3][78] = 0;
        pixel_data[3][79] = 0;
        pixel_data[3][80] = 0;
        pixel_data[3][81] = 0;
        pixel_data[3][82] = 0;
        pixel_data[3][83] = 0;
        pixel_data[3][84] = 0;
        pixel_data[3][85] = 0;
        pixel_data[3][86] = 0;
        pixel_data[3][87] = 0;
        pixel_data[3][88] = 0;
        pixel_data[3][89] = 0;
        pixel_data[3][90] = 0;
        pixel_data[3][91] = 0;
        pixel_data[3][92] = 0;
        pixel_data[3][93] = 0;
        pixel_data[3][94] = 0;
        pixel_data[3][95] = 0;
        pixel_data[3][96] = 0;
        pixel_data[3][97] = 0;
        pixel_data[3][98] = 0;
        pixel_data[3][99] = 0;
        pixel_data[3][100] = 0;
        pixel_data[3][101] = 0;
        pixel_data[3][102] = 0;
        pixel_data[3][103] = 0;
        pixel_data[3][104] = 0;
        pixel_data[3][105] = 0;
        pixel_data[3][106] = 0;
        pixel_data[3][107] = 0;
        pixel_data[3][108] = 0;
        pixel_data[3][109] = 0;
        pixel_data[3][110] = 0;
        pixel_data[3][111] = 0;
        pixel_data[3][112] = 0;
        pixel_data[3][113] = 0;
        pixel_data[3][114] = 0;
        pixel_data[3][115] = 0;
        pixel_data[3][116] = 0;
        pixel_data[3][117] = 0;
        pixel_data[3][118] = 0;
        pixel_data[3][119] = 0;
        pixel_data[3][120] = 0;
        pixel_data[3][121] = 0;
        pixel_data[3][122] = 0;
        pixel_data[3][123] = 0;
        pixel_data[3][124] = 0;
        pixel_data[3][125] = 0;
        pixel_data[3][126] = 0;
        pixel_data[3][127] = 0;
        pixel_data[3][128] = 0;
        pixel_data[3][129] = 0;
        pixel_data[3][130] = 0;
        pixel_data[3][131] = 0;
        pixel_data[3][132] = 0;
        pixel_data[3][133] = 0;
        pixel_data[3][134] = 0;
        pixel_data[3][135] = 0;
        pixel_data[3][136] = 0;
        pixel_data[3][137] = 0;
        pixel_data[3][138] = 0;
        pixel_data[3][139] = 0;
        pixel_data[3][140] = 0;
        pixel_data[3][141] = 0;
        pixel_data[3][142] = 0;
        pixel_data[3][143] = 0;
        pixel_data[3][144] = 0;
        pixel_data[3][145] = 0;
        pixel_data[3][146] = 0;
        pixel_data[3][147] = 0;
        pixel_data[3][148] = 0;
        pixel_data[3][149] = 0;
        pixel_data[3][150] = 0;
        pixel_data[3][151] = 0;
        pixel_data[3][152] = 0;
        pixel_data[3][153] = 0;
        pixel_data[3][154] = 0;
        pixel_data[3][155] = 0;
        pixel_data[3][156] = 0;
        pixel_data[3][157] = 0;
        pixel_data[3][158] = 0;
        pixel_data[3][159] = 0;
        pixel_data[3][160] = 0;
        pixel_data[3][161] = 0;
        pixel_data[3][162] = 0;
        pixel_data[3][163] = 0;
        pixel_data[3][164] = 0;
        pixel_data[3][165] = 0;
        pixel_data[3][166] = 0;
        pixel_data[3][167] = 0;
        pixel_data[3][168] = 0;
        pixel_data[3][169] = 0;
        pixel_data[3][170] = 0;
        pixel_data[3][171] = 0;
        pixel_data[3][172] = 0;
        pixel_data[3][173] = 0;
        pixel_data[3][174] = 0;
        pixel_data[3][175] = 0;
        pixel_data[3][176] = 0;
        pixel_data[3][177] = 0;
        pixel_data[3][178] = 0;
        pixel_data[3][179] = 0;
        pixel_data[3][180] = 0;
        pixel_data[3][181] = 0;
        pixel_data[3][182] = 0;
        pixel_data[3][183] = 0;
        pixel_data[3][184] = 0;
        pixel_data[3][185] = 0;
        pixel_data[3][186] = 0;
        pixel_data[3][187] = 0;
        pixel_data[3][188] = 0;
        pixel_data[3][189] = 0;
        pixel_data[3][190] = 0;
        pixel_data[3][191] = 0;
        pixel_data[3][192] = 0;
        pixel_data[3][193] = 0;
        pixel_data[3][194] = 0;
        pixel_data[3][195] = 0;
        pixel_data[3][196] = 0;
        pixel_data[3][197] = 0;
        pixel_data[3][198] = 0;
        pixel_data[3][199] = 0; // y=3
        pixel_data[4][0] = 0;
        pixel_data[4][1] = 0;
        pixel_data[4][2] = 0;
        pixel_data[4][3] = 0;
        pixel_data[4][4] = 0;
        pixel_data[4][5] = 0;
        pixel_data[4][6] = 0;
        pixel_data[4][7] = 0;
        pixel_data[4][8] = 0;
        pixel_data[4][9] = 0;
        pixel_data[4][10] = 0;
        pixel_data[4][11] = 0;
        pixel_data[4][12] = 0;
        pixel_data[4][13] = 0;
        pixel_data[4][14] = 0;
        pixel_data[4][15] = 0;
        pixel_data[4][16] = 0;
        pixel_data[4][17] = 0;
        pixel_data[4][18] = 0;
        pixel_data[4][19] = 0;
        pixel_data[4][20] = 0;
        pixel_data[4][21] = 0;
        pixel_data[4][22] = 0;
        pixel_data[4][23] = 0;
        pixel_data[4][24] = 0;
        pixel_data[4][25] = 0;
        pixel_data[4][26] = 0;
        pixel_data[4][27] = 0;
        pixel_data[4][28] = 0;
        pixel_data[4][29] = 0;
        pixel_data[4][30] = 0;
        pixel_data[4][31] = 0;
        pixel_data[4][32] = 0;
        pixel_data[4][33] = 0;
        pixel_data[4][34] = 0;
        pixel_data[4][35] = 0;
        pixel_data[4][36] = 0;
        pixel_data[4][37] = 0;
        pixel_data[4][38] = 0;
        pixel_data[4][39] = 0;
        pixel_data[4][40] = 0;
        pixel_data[4][41] = 0;
        pixel_data[4][42] = 0;
        pixel_data[4][43] = 0;
        pixel_data[4][44] = 0;
        pixel_data[4][45] = 0;
        pixel_data[4][46] = 0;
        pixel_data[4][47] = 0;
        pixel_data[4][48] = 0;
        pixel_data[4][49] = 0;
        pixel_data[4][50] = 0;
        pixel_data[4][51] = 0;
        pixel_data[4][52] = 0;
        pixel_data[4][53] = 0;
        pixel_data[4][54] = 0;
        pixel_data[4][55] = 0;
        pixel_data[4][56] = 0;
        pixel_data[4][57] = 0;
        pixel_data[4][58] = 0;
        pixel_data[4][59] = 0;
        pixel_data[4][60] = 0;
        pixel_data[4][61] = 0;
        pixel_data[4][62] = 0;
        pixel_data[4][63] = 0;
        pixel_data[4][64] = 0;
        pixel_data[4][65] = 0;
        pixel_data[4][66] = 0;
        pixel_data[4][67] = 0;
        pixel_data[4][68] = 0;
        pixel_data[4][69] = 0;
        pixel_data[4][70] = 0;
        pixel_data[4][71] = 0;
        pixel_data[4][72] = 0;
        pixel_data[4][73] = 0;
        pixel_data[4][74] = 0;
        pixel_data[4][75] = 0;
        pixel_data[4][76] = 0;
        pixel_data[4][77] = 0;
        pixel_data[4][78] = 0;
        pixel_data[4][79] = 0;
        pixel_data[4][80] = 0;
        pixel_data[4][81] = 0;
        pixel_data[4][82] = 0;
        pixel_data[4][83] = 0;
        pixel_data[4][84] = 0;
        pixel_data[4][85] = 0;
        pixel_data[4][86] = 0;
        pixel_data[4][87] = 0;
        pixel_data[4][88] = 0;
        pixel_data[4][89] = 0;
        pixel_data[4][90] = 0;
        pixel_data[4][91] = 0;
        pixel_data[4][92] = 0;
        pixel_data[4][93] = 0;
        pixel_data[4][94] = 0;
        pixel_data[4][95] = 0;
        pixel_data[4][96] = 0;
        pixel_data[4][97] = 0;
        pixel_data[4][98] = 0;
        pixel_data[4][99] = 0;
        pixel_data[4][100] = 0;
        pixel_data[4][101] = 0;
        pixel_data[4][102] = 0;
        pixel_data[4][103] = 0;
        pixel_data[4][104] = 0;
        pixel_data[4][105] = 0;
        pixel_data[4][106] = 0;
        pixel_data[4][107] = 0;
        pixel_data[4][108] = 0;
        pixel_data[4][109] = 0;
        pixel_data[4][110] = 0;
        pixel_data[4][111] = 0;
        pixel_data[4][112] = 0;
        pixel_data[4][113] = 0;
        pixel_data[4][114] = 0;
        pixel_data[4][115] = 0;
        pixel_data[4][116] = 0;
        pixel_data[4][117] = 0;
        pixel_data[4][118] = 0;
        pixel_data[4][119] = 0;
        pixel_data[4][120] = 0;
        pixel_data[4][121] = 0;
        pixel_data[4][122] = 0;
        pixel_data[4][123] = 0;
        pixel_data[4][124] = 0;
        pixel_data[4][125] = 0;
        pixel_data[4][126] = 0;
        pixel_data[4][127] = 0;
        pixel_data[4][128] = 0;
        pixel_data[4][129] = 0;
        pixel_data[4][130] = 0;
        pixel_data[4][131] = 0;
        pixel_data[4][132] = 0;
        pixel_data[4][133] = 0;
        pixel_data[4][134] = 0;
        pixel_data[4][135] = 0;
        pixel_data[4][136] = 0;
        pixel_data[4][137] = 0;
        pixel_data[4][138] = 0;
        pixel_data[4][139] = 0;
        pixel_data[4][140] = 0;
        pixel_data[4][141] = 0;
        pixel_data[4][142] = 0;
        pixel_data[4][143] = 0;
        pixel_data[4][144] = 0;
        pixel_data[4][145] = 0;
        pixel_data[4][146] = 0;
        pixel_data[4][147] = 0;
        pixel_data[4][148] = 0;
        pixel_data[4][149] = 0;
        pixel_data[4][150] = 0;
        pixel_data[4][151] = 0;
        pixel_data[4][152] = 0;
        pixel_data[4][153] = 0;
        pixel_data[4][154] = 0;
        pixel_data[4][155] = 0;
        pixel_data[4][156] = 0;
        pixel_data[4][157] = 0;
        pixel_data[4][158] = 0;
        pixel_data[4][159] = 0;
        pixel_data[4][160] = 0;
        pixel_data[4][161] = 0;
        pixel_data[4][162] = 0;
        pixel_data[4][163] = 0;
        pixel_data[4][164] = 0;
        pixel_data[4][165] = 0;
        pixel_data[4][166] = 0;
        pixel_data[4][167] = 0;
        pixel_data[4][168] = 0;
        pixel_data[4][169] = 0;
        pixel_data[4][170] = 0;
        pixel_data[4][171] = 0;
        pixel_data[4][172] = 0;
        pixel_data[4][173] = 0;
        pixel_data[4][174] = 0;
        pixel_data[4][175] = 0;
        pixel_data[4][176] = 0;
        pixel_data[4][177] = 0;
        pixel_data[4][178] = 0;
        pixel_data[4][179] = 0;
        pixel_data[4][180] = 0;
        pixel_data[4][181] = 0;
        pixel_data[4][182] = 0;
        pixel_data[4][183] = 0;
        pixel_data[4][184] = 0;
        pixel_data[4][185] = 0;
        pixel_data[4][186] = 0;
        pixel_data[4][187] = 0;
        pixel_data[4][188] = 0;
        pixel_data[4][189] = 0;
        pixel_data[4][190] = 0;
        pixel_data[4][191] = 0;
        pixel_data[4][192] = 0;
        pixel_data[4][193] = 0;
        pixel_data[4][194] = 0;
        pixel_data[4][195] = 0;
        pixel_data[4][196] = 0;
        pixel_data[4][197] = 0;
        pixel_data[4][198] = 0;
        pixel_data[4][199] = 0; // y=4
        pixel_data[5][0] = 0;
        pixel_data[5][1] = 0;
        pixel_data[5][2] = 0;
        pixel_data[5][3] = 0;
        pixel_data[5][4] = 0;
        pixel_data[5][5] = 0;
        pixel_data[5][6] = 0;
        pixel_data[5][7] = 0;
        pixel_data[5][8] = 0;
        pixel_data[5][9] = 0;
        pixel_data[5][10] = 0;
        pixel_data[5][11] = 0;
        pixel_data[5][12] = 0;
        pixel_data[5][13] = 0;
        pixel_data[5][14] = 0;
        pixel_data[5][15] = 0;
        pixel_data[5][16] = 0;
        pixel_data[5][17] = 0;
        pixel_data[5][18] = 0;
        pixel_data[5][19] = 0;
        pixel_data[5][20] = 0;
        pixel_data[5][21] = 0;
        pixel_data[5][22] = 0;
        pixel_data[5][23] = 0;
        pixel_data[5][24] = 0;
        pixel_data[5][25] = 0;
        pixel_data[5][26] = 0;
        pixel_data[5][27] = 0;
        pixel_data[5][28] = 0;
        pixel_data[5][29] = 0;
        pixel_data[5][30] = 0;
        pixel_data[5][31] = 0;
        pixel_data[5][32] = 0;
        pixel_data[5][33] = 0;
        pixel_data[5][34] = 0;
        pixel_data[5][35] = 0;
        pixel_data[5][36] = 0;
        pixel_data[5][37] = 0;
        pixel_data[5][38] = 0;
        pixel_data[5][39] = 0;
        pixel_data[5][40] = 0;
        pixel_data[5][41] = 0;
        pixel_data[5][42] = 0;
        pixel_data[5][43] = 0;
        pixel_data[5][44] = 0;
        pixel_data[5][45] = 0;
        pixel_data[5][46] = 0;
        pixel_data[5][47] = 0;
        pixel_data[5][48] = 0;
        pixel_data[5][49] = 0;
        pixel_data[5][50] = 0;
        pixel_data[5][51] = 0;
        pixel_data[5][52] = 0;
        pixel_data[5][53] = 0;
        pixel_data[5][54] = 0;
        pixel_data[5][55] = 0;
        pixel_data[5][56] = 0;
        pixel_data[5][57] = 0;
        pixel_data[5][58] = 0;
        pixel_data[5][59] = 0;
        pixel_data[5][60] = 0;
        pixel_data[5][61] = 0;
        pixel_data[5][62] = 0;
        pixel_data[5][63] = 0;
        pixel_data[5][64] = 0;
        pixel_data[5][65] = 0;
        pixel_data[5][66] = 0;
        pixel_data[5][67] = 0;
        pixel_data[5][68] = 0;
        pixel_data[5][69] = 0;
        pixel_data[5][70] = 0;
        pixel_data[5][71] = 0;
        pixel_data[5][72] = 0;
        pixel_data[5][73] = 0;
        pixel_data[5][74] = 0;
        pixel_data[5][75] = 0;
        pixel_data[5][76] = 0;
        pixel_data[5][77] = 0;
        pixel_data[5][78] = 0;
        pixel_data[5][79] = 0;
        pixel_data[5][80] = 0;
        pixel_data[5][81] = 0;
        pixel_data[5][82] = 0;
        pixel_data[5][83] = 0;
        pixel_data[5][84] = 0;
        pixel_data[5][85] = 0;
        pixel_data[5][86] = 0;
        pixel_data[5][87] = 0;
        pixel_data[5][88] = 0;
        pixel_data[5][89] = 0;
        pixel_data[5][90] = 0;
        pixel_data[5][91] = 0;
        pixel_data[5][92] = 0;
        pixel_data[5][93] = 0;
        pixel_data[5][94] = 0;
        pixel_data[5][95] = 0;
        pixel_data[5][96] = 0;
        pixel_data[5][97] = 0;
        pixel_data[5][98] = 0;
        pixel_data[5][99] = 0;
        pixel_data[5][100] = 0;
        pixel_data[5][101] = 0;
        pixel_data[5][102] = 0;
        pixel_data[5][103] = 0;
        pixel_data[5][104] = 0;
        pixel_data[5][105] = 0;
        pixel_data[5][106] = 0;
        pixel_data[5][107] = 0;
        pixel_data[5][108] = 0;
        pixel_data[5][109] = 0;
        pixel_data[5][110] = 0;
        pixel_data[5][111] = 0;
        pixel_data[5][112] = 0;
        pixel_data[5][113] = 0;
        pixel_data[5][114] = 0;
        pixel_data[5][115] = 0;
        pixel_data[5][116] = 0;
        pixel_data[5][117] = 0;
        pixel_data[5][118] = 0;
        pixel_data[5][119] = 0;
        pixel_data[5][120] = 0;
        pixel_data[5][121] = 0;
        pixel_data[5][122] = 0;
        pixel_data[5][123] = 0;
        pixel_data[5][124] = 0;
        pixel_data[5][125] = 0;
        pixel_data[5][126] = 0;
        pixel_data[5][127] = 0;
        pixel_data[5][128] = 0;
        pixel_data[5][129] = 0;
        pixel_data[5][130] = 0;
        pixel_data[5][131] = 0;
        pixel_data[5][132] = 0;
        pixel_data[5][133] = 0;
        pixel_data[5][134] = 0;
        pixel_data[5][135] = 0;
        pixel_data[5][136] = 0;
        pixel_data[5][137] = 0;
        pixel_data[5][138] = 0;
        pixel_data[5][139] = 0;
        pixel_data[5][140] = 0;
        pixel_data[5][141] = 0;
        pixel_data[5][142] = 0;
        pixel_data[5][143] = 0;
        pixel_data[5][144] = 0;
        pixel_data[5][145] = 0;
        pixel_data[5][146] = 0;
        pixel_data[5][147] = 0;
        pixel_data[5][148] = 0;
        pixel_data[5][149] = 0;
        pixel_data[5][150] = 0;
        pixel_data[5][151] = 0;
        pixel_data[5][152] = 0;
        pixel_data[5][153] = 0;
        pixel_data[5][154] = 0;
        pixel_data[5][155] = 0;
        pixel_data[5][156] = 0;
        pixel_data[5][157] = 0;
        pixel_data[5][158] = 0;
        pixel_data[5][159] = 0;
        pixel_data[5][160] = 0;
        pixel_data[5][161] = 0;
        pixel_data[5][162] = 0;
        pixel_data[5][163] = 0;
        pixel_data[5][164] = 0;
        pixel_data[5][165] = 0;
        pixel_data[5][166] = 0;
        pixel_data[5][167] = 0;
        pixel_data[5][168] = 0;
        pixel_data[5][169] = 0;
        pixel_data[5][170] = 0;
        pixel_data[5][171] = 0;
        pixel_data[5][172] = 0;
        pixel_data[5][173] = 0;
        pixel_data[5][174] = 0;
        pixel_data[5][175] = 0;
        pixel_data[5][176] = 0;
        pixel_data[5][177] = 0;
        pixel_data[5][178] = 0;
        pixel_data[5][179] = 0;
        pixel_data[5][180] = 0;
        pixel_data[5][181] = 0;
        pixel_data[5][182] = 0;
        pixel_data[5][183] = 0;
        pixel_data[5][184] = 0;
        pixel_data[5][185] = 0;
        pixel_data[5][186] = 0;
        pixel_data[5][187] = 0;
        pixel_data[5][188] = 0;
        pixel_data[5][189] = 0;
        pixel_data[5][190] = 0;
        pixel_data[5][191] = 0;
        pixel_data[5][192] = 0;
        pixel_data[5][193] = 0;
        pixel_data[5][194] = 0;
        pixel_data[5][195] = 0;
        pixel_data[5][196] = 0;
        pixel_data[5][197] = 0;
        pixel_data[5][198] = 0;
        pixel_data[5][199] = 0; // y=5
        pixel_data[6][0] = 0;
        pixel_data[6][1] = 0;
        pixel_data[6][2] = 0;
        pixel_data[6][3] = 0;
        pixel_data[6][4] = 0;
        pixel_data[6][5] = 0;
        pixel_data[6][6] = 0;
        pixel_data[6][7] = 0;
        pixel_data[6][8] = 0;
        pixel_data[6][9] = 0;
        pixel_data[6][10] = 0;
        pixel_data[6][11] = 0;
        pixel_data[6][12] = 0;
        pixel_data[6][13] = 0;
        pixel_data[6][14] = 0;
        pixel_data[6][15] = 0;
        pixel_data[6][16] = 0;
        pixel_data[6][17] = 0;
        pixel_data[6][18] = 0;
        pixel_data[6][19] = 0;
        pixel_data[6][20] = 0;
        pixel_data[6][21] = 0;
        pixel_data[6][22] = 0;
        pixel_data[6][23] = 0;
        pixel_data[6][24] = 0;
        pixel_data[6][25] = 0;
        pixel_data[6][26] = 0;
        pixel_data[6][27] = 0;
        pixel_data[6][28] = 0;
        pixel_data[6][29] = 0;
        pixel_data[6][30] = 0;
        pixel_data[6][31] = 0;
        pixel_data[6][32] = 0;
        pixel_data[6][33] = 0;
        pixel_data[6][34] = 0;
        pixel_data[6][35] = 0;
        pixel_data[6][36] = 0;
        pixel_data[6][37] = 0;
        pixel_data[6][38] = 0;
        pixel_data[6][39] = 0;
        pixel_data[6][40] = 0;
        pixel_data[6][41] = 0;
        pixel_data[6][42] = 0;
        pixel_data[6][43] = 0;
        pixel_data[6][44] = 0;
        pixel_data[6][45] = 0;
        pixel_data[6][46] = 0;
        pixel_data[6][47] = 0;
        pixel_data[6][48] = 0;
        pixel_data[6][49] = 0;
        pixel_data[6][50] = 0;
        pixel_data[6][51] = 0;
        pixel_data[6][52] = 0;
        pixel_data[6][53] = 0;
        pixel_data[6][54] = 0;
        pixel_data[6][55] = 0;
        pixel_data[6][56] = 0;
        pixel_data[6][57] = 0;
        pixel_data[6][58] = 0;
        pixel_data[6][59] = 0;
        pixel_data[6][60] = 0;
        pixel_data[6][61] = 0;
        pixel_data[6][62] = 0;
        pixel_data[6][63] = 0;
        pixel_data[6][64] = 0;
        pixel_data[6][65] = 0;
        pixel_data[6][66] = 0;
        pixel_data[6][67] = 0;
        pixel_data[6][68] = 0;
        pixel_data[6][69] = 0;
        pixel_data[6][70] = 0;
        pixel_data[6][71] = 0;
        pixel_data[6][72] = 0;
        pixel_data[6][73] = 0;
        pixel_data[6][74] = 0;
        pixel_data[6][75] = 0;
        pixel_data[6][76] = 0;
        pixel_data[6][77] = 0;
        pixel_data[6][78] = 0;
        pixel_data[6][79] = 0;
        pixel_data[6][80] = 0;
        pixel_data[6][81] = 0;
        pixel_data[6][82] = 0;
        pixel_data[6][83] = 0;
        pixel_data[6][84] = 0;
        pixel_data[6][85] = 0;
        pixel_data[6][86] = 0;
        pixel_data[6][87] = 0;
        pixel_data[6][88] = 0;
        pixel_data[6][89] = 0;
        pixel_data[6][90] = 0;
        pixel_data[6][91] = 0;
        pixel_data[6][92] = 0;
        pixel_data[6][93] = 0;
        pixel_data[6][94] = 0;
        pixel_data[6][95] = 0;
        pixel_data[6][96] = 0;
        pixel_data[6][97] = 0;
        pixel_data[6][98] = 0;
        pixel_data[6][99] = 0;
        pixel_data[6][100] = 0;
        pixel_data[6][101] = 0;
        pixel_data[6][102] = 0;
        pixel_data[6][103] = 0;
        pixel_data[6][104] = 0;
        pixel_data[6][105] = 0;
        pixel_data[6][106] = 0;
        pixel_data[6][107] = 0;
        pixel_data[6][108] = 0;
        pixel_data[6][109] = 0;
        pixel_data[6][110] = 0;
        pixel_data[6][111] = 0;
        pixel_data[6][112] = 0;
        pixel_data[6][113] = 0;
        pixel_data[6][114] = 0;
        pixel_data[6][115] = 0;
        pixel_data[6][116] = 0;
        pixel_data[6][117] = 0;
        pixel_data[6][118] = 0;
        pixel_data[6][119] = 0;
        pixel_data[6][120] = 0;
        pixel_data[6][121] = 0;
        pixel_data[6][122] = 0;
        pixel_data[6][123] = 0;
        pixel_data[6][124] = 0;
        pixel_data[6][125] = 0;
        pixel_data[6][126] = 0;
        pixel_data[6][127] = 0;
        pixel_data[6][128] = 0;
        pixel_data[6][129] = 0;
        pixel_data[6][130] = 0;
        pixel_data[6][131] = 0;
        pixel_data[6][132] = 0;
        pixel_data[6][133] = 0;
        pixel_data[6][134] = 0;
        pixel_data[6][135] = 0;
        pixel_data[6][136] = 0;
        pixel_data[6][137] = 0;
        pixel_data[6][138] = 0;
        pixel_data[6][139] = 0;
        pixel_data[6][140] = 0;
        pixel_data[6][141] = 0;
        pixel_data[6][142] = 0;
        pixel_data[6][143] = 0;
        pixel_data[6][144] = 0;
        pixel_data[6][145] = 0;
        pixel_data[6][146] = 0;
        pixel_data[6][147] = 0;
        pixel_data[6][148] = 0;
        pixel_data[6][149] = 0;
        pixel_data[6][150] = 0;
        pixel_data[6][151] = 0;
        pixel_data[6][152] = 0;
        pixel_data[6][153] = 0;
        pixel_data[6][154] = 0;
        pixel_data[6][155] = 0;
        pixel_data[6][156] = 0;
        pixel_data[6][157] = 0;
        pixel_data[6][158] = 0;
        pixel_data[6][159] = 0;
        pixel_data[6][160] = 0;
        pixel_data[6][161] = 0;
        pixel_data[6][162] = 0;
        pixel_data[6][163] = 0;
        pixel_data[6][164] = 0;
        pixel_data[6][165] = 0;
        pixel_data[6][166] = 0;
        pixel_data[6][167] = 0;
        pixel_data[6][168] = 0;
        pixel_data[6][169] = 0;
        pixel_data[6][170] = 0;
        pixel_data[6][171] = 0;
        pixel_data[6][172] = 0;
        pixel_data[6][173] = 0;
        pixel_data[6][174] = 0;
        pixel_data[6][175] = 0;
        pixel_data[6][176] = 0;
        pixel_data[6][177] = 0;
        pixel_data[6][178] = 0;
        pixel_data[6][179] = 0;
        pixel_data[6][180] = 0;
        pixel_data[6][181] = 0;
        pixel_data[6][182] = 0;
        pixel_data[6][183] = 0;
        pixel_data[6][184] = 0;
        pixel_data[6][185] = 0;
        pixel_data[6][186] = 0;
        pixel_data[6][187] = 0;
        pixel_data[6][188] = 0;
        pixel_data[6][189] = 0;
        pixel_data[6][190] = 0;
        pixel_data[6][191] = 0;
        pixel_data[6][192] = 0;
        pixel_data[6][193] = 0;
        pixel_data[6][194] = 0;
        pixel_data[6][195] = 0;
        pixel_data[6][196] = 0;
        pixel_data[6][197] = 0;
        pixel_data[6][198] = 0;
        pixel_data[6][199] = 0; // y=6
        pixel_data[7][0] = 0;
        pixel_data[7][1] = 0;
        pixel_data[7][2] = 0;
        pixel_data[7][3] = 0;
        pixel_data[7][4] = 0;
        pixel_data[7][5] = 0;
        pixel_data[7][6] = 0;
        pixel_data[7][7] = 0;
        pixel_data[7][8] = 0;
        pixel_data[7][9] = 0;
        pixel_data[7][10] = 0;
        pixel_data[7][11] = 0;
        pixel_data[7][12] = 0;
        pixel_data[7][13] = 0;
        pixel_data[7][14] = 0;
        pixel_data[7][15] = 0;
        pixel_data[7][16] = 0;
        pixel_data[7][17] = 0;
        pixel_data[7][18] = 0;
        pixel_data[7][19] = 0;
        pixel_data[7][20] = 0;
        pixel_data[7][21] = 0;
        pixel_data[7][22] = 0;
        pixel_data[7][23] = 0;
        pixel_data[7][24] = 0;
        pixel_data[7][25] = 0;
        pixel_data[7][26] = 0;
        pixel_data[7][27] = 0;
        pixel_data[7][28] = 0;
        pixel_data[7][29] = 0;
        pixel_data[7][30] = 0;
        pixel_data[7][31] = 0;
        pixel_data[7][32] = 0;
        pixel_data[7][33] = 0;
        pixel_data[7][34] = 0;
        pixel_data[7][35] = 0;
        pixel_data[7][36] = 0;
        pixel_data[7][37] = 0;
        pixel_data[7][38] = 0;
        pixel_data[7][39] = 0;
        pixel_data[7][40] = 0;
        pixel_data[7][41] = 0;
        pixel_data[7][42] = 0;
        pixel_data[7][43] = 0;
        pixel_data[7][44] = 0;
        pixel_data[7][45] = 0;
        pixel_data[7][46] = 0;
        pixel_data[7][47] = 0;
        pixel_data[7][48] = 0;
        pixel_data[7][49] = 0;
        pixel_data[7][50] = 0;
        pixel_data[7][51] = 0;
        pixel_data[7][52] = 0;
        pixel_data[7][53] = 0;
        pixel_data[7][54] = 0;
        pixel_data[7][55] = 0;
        pixel_data[7][56] = 0;
        pixel_data[7][57] = 0;
        pixel_data[7][58] = 0;
        pixel_data[7][59] = 0;
        pixel_data[7][60] = 0;
        pixel_data[7][61] = 0;
        pixel_data[7][62] = 0;
        pixel_data[7][63] = 0;
        pixel_data[7][64] = 0;
        pixel_data[7][65] = 0;
        pixel_data[7][66] = 0;
        pixel_data[7][67] = 0;
        pixel_data[7][68] = 0;
        pixel_data[7][69] = 0;
        pixel_data[7][70] = 0;
        pixel_data[7][71] = 0;
        pixel_data[7][72] = 0;
        pixel_data[7][73] = 0;
        pixel_data[7][74] = 0;
        pixel_data[7][75] = 0;
        pixel_data[7][76] = 0;
        pixel_data[7][77] = 0;
        pixel_data[7][78] = 0;
        pixel_data[7][79] = 0;
        pixel_data[7][80] = 0;
        pixel_data[7][81] = 0;
        pixel_data[7][82] = 0;
        pixel_data[7][83] = 0;
        pixel_data[7][84] = 0;
        pixel_data[7][85] = 0;
        pixel_data[7][86] = 0;
        pixel_data[7][87] = 0;
        pixel_data[7][88] = 0;
        pixel_data[7][89] = 0;
        pixel_data[7][90] = 0;
        pixel_data[7][91] = 0;
        pixel_data[7][92] = 0;
        pixel_data[7][93] = 0;
        pixel_data[7][94] = 0;
        pixel_data[7][95] = 0;
        pixel_data[7][96] = 0;
        pixel_data[7][97] = 0;
        pixel_data[7][98] = 0;
        pixel_data[7][99] = 0;
        pixel_data[7][100] = 0;
        pixel_data[7][101] = 0;
        pixel_data[7][102] = 0;
        pixel_data[7][103] = 0;
        pixel_data[7][104] = 0;
        pixel_data[7][105] = 0;
        pixel_data[7][106] = 0;
        pixel_data[7][107] = 0;
        pixel_data[7][108] = 0;
        pixel_data[7][109] = 0;
        pixel_data[7][110] = 0;
        pixel_data[7][111] = 0;
        pixel_data[7][112] = 0;
        pixel_data[7][113] = 0;
        pixel_data[7][114] = 0;
        pixel_data[7][115] = 0;
        pixel_data[7][116] = 0;
        pixel_data[7][117] = 0;
        pixel_data[7][118] = 0;
        pixel_data[7][119] = 0;
        pixel_data[7][120] = 0;
        pixel_data[7][121] = 0;
        pixel_data[7][122] = 0;
        pixel_data[7][123] = 0;
        pixel_data[7][124] = 0;
        pixel_data[7][125] = 0;
        pixel_data[7][126] = 0;
        pixel_data[7][127] = 0;
        pixel_data[7][128] = 0;
        pixel_data[7][129] = 0;
        pixel_data[7][130] = 0;
        pixel_data[7][131] = 0;
        pixel_data[7][132] = 0;
        pixel_data[7][133] = 0;
        pixel_data[7][134] = 0;
        pixel_data[7][135] = 0;
        pixel_data[7][136] = 0;
        pixel_data[7][137] = 0;
        pixel_data[7][138] = 0;
        pixel_data[7][139] = 0;
        pixel_data[7][140] = 0;
        pixel_data[7][141] = 0;
        pixel_data[7][142] = 0;
        pixel_data[7][143] = 0;
        pixel_data[7][144] = 0;
        pixel_data[7][145] = 0;
        pixel_data[7][146] = 0;
        pixel_data[7][147] = 0;
        pixel_data[7][148] = 0;
        pixel_data[7][149] = 0;
        pixel_data[7][150] = 0;
        pixel_data[7][151] = 0;
        pixel_data[7][152] = 0;
        pixel_data[7][153] = 0;
        pixel_data[7][154] = 0;
        pixel_data[7][155] = 0;
        pixel_data[7][156] = 0;
        pixel_data[7][157] = 0;
        pixel_data[7][158] = 0;
        pixel_data[7][159] = 0;
        pixel_data[7][160] = 0;
        pixel_data[7][161] = 0;
        pixel_data[7][162] = 0;
        pixel_data[7][163] = 0;
        pixel_data[7][164] = 0;
        pixel_data[7][165] = 0;
        pixel_data[7][166] = 0;
        pixel_data[7][167] = 0;
        pixel_data[7][168] = 0;
        pixel_data[7][169] = 0;
        pixel_data[7][170] = 0;
        pixel_data[7][171] = 0;
        pixel_data[7][172] = 0;
        pixel_data[7][173] = 0;
        pixel_data[7][174] = 0;
        pixel_data[7][175] = 0;
        pixel_data[7][176] = 0;
        pixel_data[7][177] = 0;
        pixel_data[7][178] = 0;
        pixel_data[7][179] = 0;
        pixel_data[7][180] = 0;
        pixel_data[7][181] = 0;
        pixel_data[7][182] = 0;
        pixel_data[7][183] = 0;
        pixel_data[7][184] = 0;
        pixel_data[7][185] = 0;
        pixel_data[7][186] = 0;
        pixel_data[7][187] = 0;
        pixel_data[7][188] = 0;
        pixel_data[7][189] = 0;
        pixel_data[7][190] = 0;
        pixel_data[7][191] = 0;
        pixel_data[7][192] = 0;
        pixel_data[7][193] = 0;
        pixel_data[7][194] = 0;
        pixel_data[7][195] = 0;
        pixel_data[7][196] = 0;
        pixel_data[7][197] = 0;
        pixel_data[7][198] = 0;
        pixel_data[7][199] = 0; // y=7
        pixel_data[8][0] = 0;
        pixel_data[8][1] = 0;
        pixel_data[8][2] = 0;
        pixel_data[8][3] = 0;
        pixel_data[8][4] = 0;
        pixel_data[8][5] = 0;
        pixel_data[8][6] = 0;
        pixel_data[8][7] = 0;
        pixel_data[8][8] = 0;
        pixel_data[8][9] = 0;
        pixel_data[8][10] = 0;
        pixel_data[8][11] = 0;
        pixel_data[8][12] = 0;
        pixel_data[8][13] = 0;
        pixel_data[8][14] = 0;
        pixel_data[8][15] = 0;
        pixel_data[8][16] = 0;
        pixel_data[8][17] = 0;
        pixel_data[8][18] = 0;
        pixel_data[8][19] = 0;
        pixel_data[8][20] = 0;
        pixel_data[8][21] = 0;
        pixel_data[8][22] = 0;
        pixel_data[8][23] = 0;
        pixel_data[8][24] = 0;
        pixel_data[8][25] = 0;
        pixel_data[8][26] = 0;
        pixel_data[8][27] = 0;
        pixel_data[8][28] = 0;
        pixel_data[8][29] = 0;
        pixel_data[8][30] = 0;
        pixel_data[8][31] = 0;
        pixel_data[8][32] = 0;
        pixel_data[8][33] = 0;
        pixel_data[8][34] = 0;
        pixel_data[8][35] = 0;
        pixel_data[8][36] = 0;
        pixel_data[8][37] = 0;
        pixel_data[8][38] = 0;
        pixel_data[8][39] = 0;
        pixel_data[8][40] = 0;
        pixel_data[8][41] = 0;
        pixel_data[8][42] = 0;
        pixel_data[8][43] = 0;
        pixel_data[8][44] = 0;
        pixel_data[8][45] = 0;
        pixel_data[8][46] = 0;
        pixel_data[8][47] = 0;
        pixel_data[8][48] = 0;
        pixel_data[8][49] = 0;
        pixel_data[8][50] = 0;
        pixel_data[8][51] = 0;
        pixel_data[8][52] = 0;
        pixel_data[8][53] = 0;
        pixel_data[8][54] = 0;
        pixel_data[8][55] = 0;
        pixel_data[8][56] = 0;
        pixel_data[8][57] = 0;
        pixel_data[8][58] = 0;
        pixel_data[8][59] = 0;
        pixel_data[8][60] = 0;
        pixel_data[8][61] = 0;
        pixel_data[8][62] = 0;
        pixel_data[8][63] = 0;
        pixel_data[8][64] = 0;
        pixel_data[8][65] = 0;
        pixel_data[8][66] = 0;
        pixel_data[8][67] = 0;
        pixel_data[8][68] = 0;
        pixel_data[8][69] = 0;
        pixel_data[8][70] = 0;
        pixel_data[8][71] = 0;
        pixel_data[8][72] = 0;
        pixel_data[8][73] = 0;
        pixel_data[8][74] = 0;
        pixel_data[8][75] = 0;
        pixel_data[8][76] = 0;
        pixel_data[8][77] = 0;
        pixel_data[8][78] = 0;
        pixel_data[8][79] = 0;
        pixel_data[8][80] = 0;
        pixel_data[8][81] = 0;
        pixel_data[8][82] = 0;
        pixel_data[8][83] = 0;
        pixel_data[8][84] = 0;
        pixel_data[8][85] = 0;
        pixel_data[8][86] = 0;
        pixel_data[8][87] = 0;
        pixel_data[8][88] = 0;
        pixel_data[8][89] = 0;
        pixel_data[8][90] = 0;
        pixel_data[8][91] = 0;
        pixel_data[8][92] = 0;
        pixel_data[8][93] = 0;
        pixel_data[8][94] = 0;
        pixel_data[8][95] = 0;
        pixel_data[8][96] = 0;
        pixel_data[8][97] = 0;
        pixel_data[8][98] = 0;
        pixel_data[8][99] = 0;
        pixel_data[8][100] = 0;
        pixel_data[8][101] = 0;
        pixel_data[8][102] = 0;
        pixel_data[8][103] = 0;
        pixel_data[8][104] = 0;
        pixel_data[8][105] = 0;
        pixel_data[8][106] = 0;
        pixel_data[8][107] = 0;
        pixel_data[8][108] = 0;
        pixel_data[8][109] = 0;
        pixel_data[8][110] = 0;
        pixel_data[8][111] = 0;
        pixel_data[8][112] = 0;
        pixel_data[8][113] = 0;
        pixel_data[8][114] = 0;
        pixel_data[8][115] = 0;
        pixel_data[8][116] = 0;
        pixel_data[8][117] = 0;
        pixel_data[8][118] = 0;
        pixel_data[8][119] = 0;
        pixel_data[8][120] = 0;
        pixel_data[8][121] = 0;
        pixel_data[8][122] = 0;
        pixel_data[8][123] = 0;
        pixel_data[8][124] = 0;
        pixel_data[8][125] = 0;
        pixel_data[8][126] = 0;
        pixel_data[8][127] = 0;
        pixel_data[8][128] = 0;
        pixel_data[8][129] = 0;
        pixel_data[8][130] = 0;
        pixel_data[8][131] = 0;
        pixel_data[8][132] = 0;
        pixel_data[8][133] = 0;
        pixel_data[8][134] = 0;
        pixel_data[8][135] = 0;
        pixel_data[8][136] = 0;
        pixel_data[8][137] = 0;
        pixel_data[8][138] = 0;
        pixel_data[8][139] = 0;
        pixel_data[8][140] = 0;
        pixel_data[8][141] = 0;
        pixel_data[8][142] = 0;
        pixel_data[8][143] = 0;
        pixel_data[8][144] = 0;
        pixel_data[8][145] = 0;
        pixel_data[8][146] = 0;
        pixel_data[8][147] = 0;
        pixel_data[8][148] = 0;
        pixel_data[8][149] = 0;
        pixel_data[8][150] = 0;
        pixel_data[8][151] = 0;
        pixel_data[8][152] = 0;
        pixel_data[8][153] = 0;
        pixel_data[8][154] = 0;
        pixel_data[8][155] = 0;
        pixel_data[8][156] = 0;
        pixel_data[8][157] = 0;
        pixel_data[8][158] = 0;
        pixel_data[8][159] = 0;
        pixel_data[8][160] = 0;
        pixel_data[8][161] = 0;
        pixel_data[8][162] = 0;
        pixel_data[8][163] = 0;
        pixel_data[8][164] = 0;
        pixel_data[8][165] = 0;
        pixel_data[8][166] = 0;
        pixel_data[8][167] = 0;
        pixel_data[8][168] = 0;
        pixel_data[8][169] = 0;
        pixel_data[8][170] = 0;
        pixel_data[8][171] = 0;
        pixel_data[8][172] = 0;
        pixel_data[8][173] = 0;
        pixel_data[8][174] = 0;
        pixel_data[8][175] = 0;
        pixel_data[8][176] = 0;
        pixel_data[8][177] = 0;
        pixel_data[8][178] = 0;
        pixel_data[8][179] = 0;
        pixel_data[8][180] = 0;
        pixel_data[8][181] = 0;
        pixel_data[8][182] = 0;
        pixel_data[8][183] = 0;
        pixel_data[8][184] = 0;
        pixel_data[8][185] = 0;
        pixel_data[8][186] = 0;
        pixel_data[8][187] = 0;
        pixel_data[8][188] = 0;
        pixel_data[8][189] = 0;
        pixel_data[8][190] = 0;
        pixel_data[8][191] = 0;
        pixel_data[8][192] = 0;
        pixel_data[8][193] = 0;
        pixel_data[8][194] = 0;
        pixel_data[8][195] = 0;
        pixel_data[8][196] = 0;
        pixel_data[8][197] = 0;
        pixel_data[8][198] = 0;
        pixel_data[8][199] = 0; // y=8
        pixel_data[9][0] = 0;
        pixel_data[9][1] = 0;
        pixel_data[9][2] = 0;
        pixel_data[9][3] = 0;
        pixel_data[9][4] = 0;
        pixel_data[9][5] = 0;
        pixel_data[9][6] = 0;
        pixel_data[9][7] = 0;
        pixel_data[9][8] = 0;
        pixel_data[9][9] = 0;
        pixel_data[9][10] = 0;
        pixel_data[9][11] = 0;
        pixel_data[9][12] = 0;
        pixel_data[9][13] = 0;
        pixel_data[9][14] = 0;
        pixel_data[9][15] = 0;
        pixel_data[9][16] = 0;
        pixel_data[9][17] = 0;
        pixel_data[9][18] = 0;
        pixel_data[9][19] = 0;
        pixel_data[9][20] = 0;
        pixel_data[9][21] = 0;
        pixel_data[9][22] = 0;
        pixel_data[9][23] = 0;
        pixel_data[9][24] = 0;
        pixel_data[9][25] = 0;
        pixel_data[9][26] = 0;
        pixel_data[9][27] = 0;
        pixel_data[9][28] = 0;
        pixel_data[9][29] = 0;
        pixel_data[9][30] = 0;
        pixel_data[9][31] = 0;
        pixel_data[9][32] = 0;
        pixel_data[9][33] = 0;
        pixel_data[9][34] = 0;
        pixel_data[9][35] = 0;
        pixel_data[9][36] = 0;
        pixel_data[9][37] = 0;
        pixel_data[9][38] = 0;
        pixel_data[9][39] = 0;
        pixel_data[9][40] = 0;
        pixel_data[9][41] = 0;
        pixel_data[9][42] = 0;
        pixel_data[9][43] = 0;
        pixel_data[9][44] = 0;
        pixel_data[9][45] = 0;
        pixel_data[9][46] = 0;
        pixel_data[9][47] = 0;
        pixel_data[9][48] = 0;
        pixel_data[9][49] = 0;
        pixel_data[9][50] = 0;
        pixel_data[9][51] = 0;
        pixel_data[9][52] = 0;
        pixel_data[9][53] = 0;
        pixel_data[9][54] = 0;
        pixel_data[9][55] = 0;
        pixel_data[9][56] = 0;
        pixel_data[9][57] = 0;
        pixel_data[9][58] = 0;
        pixel_data[9][59] = 0;
        pixel_data[9][60] = 0;
        pixel_data[9][61] = 0;
        pixel_data[9][62] = 0;
        pixel_data[9][63] = 0;
        pixel_data[9][64] = 0;
        pixel_data[9][65] = 0;
        pixel_data[9][66] = 0;
        pixel_data[9][67] = 0;
        pixel_data[9][68] = 0;
        pixel_data[9][69] = 0;
        pixel_data[9][70] = 0;
        pixel_data[9][71] = 0;
        pixel_data[9][72] = 0;
        pixel_data[9][73] = 0;
        pixel_data[9][74] = 0;
        pixel_data[9][75] = 0;
        pixel_data[9][76] = 0;
        pixel_data[9][77] = 0;
        pixel_data[9][78] = 0;
        pixel_data[9][79] = 0;
        pixel_data[9][80] = 0;
        pixel_data[9][81] = 0;
        pixel_data[9][82] = 0;
        pixel_data[9][83] = 0;
        pixel_data[9][84] = 0;
        pixel_data[9][85] = 0;
        pixel_data[9][86] = 0;
        pixel_data[9][87] = 0;
        pixel_data[9][88] = 0;
        pixel_data[9][89] = 0;
        pixel_data[9][90] = 0;
        pixel_data[9][91] = 0;
        pixel_data[9][92] = 0;
        pixel_data[9][93] = 0;
        pixel_data[9][94] = 0;
        pixel_data[9][95] = 0;
        pixel_data[9][96] = 0;
        pixel_data[9][97] = 0;
        pixel_data[9][98] = 0;
        pixel_data[9][99] = 0;
        pixel_data[9][100] = 0;
        pixel_data[9][101] = 0;
        pixel_data[9][102] = 0;
        pixel_data[9][103] = 0;
        pixel_data[9][104] = 0;
        pixel_data[9][105] = 0;
        pixel_data[9][106] = 0;
        pixel_data[9][107] = 0;
        pixel_data[9][108] = 0;
        pixel_data[9][109] = 0;
        pixel_data[9][110] = 0;
        pixel_data[9][111] = 0;
        pixel_data[9][112] = 0;
        pixel_data[9][113] = 0;
        pixel_data[9][114] = 0;
        pixel_data[9][115] = 0;
        pixel_data[9][116] = 0;
        pixel_data[9][117] = 0;
        pixel_data[9][118] = 0;
        pixel_data[9][119] = 0;
        pixel_data[9][120] = 0;
        pixel_data[9][121] = 0;
        pixel_data[9][122] = 0;
        pixel_data[9][123] = 0;
        pixel_data[9][124] = 0;
        pixel_data[9][125] = 0;
        pixel_data[9][126] = 0;
        pixel_data[9][127] = 0;
        pixel_data[9][128] = 0;
        pixel_data[9][129] = 0;
        pixel_data[9][130] = 0;
        pixel_data[9][131] = 0;
        pixel_data[9][132] = 0;
        pixel_data[9][133] = 0;
        pixel_data[9][134] = 0;
        pixel_data[9][135] = 0;
        pixel_data[9][136] = 0;
        pixel_data[9][137] = 0;
        pixel_data[9][138] = 0;
        pixel_data[9][139] = 0;
        pixel_data[9][140] = 0;
        pixel_data[9][141] = 0;
        pixel_data[9][142] = 0;
        pixel_data[9][143] = 0;
        pixel_data[9][144] = 0;
        pixel_data[9][145] = 0;
        pixel_data[9][146] = 0;
        pixel_data[9][147] = 0;
        pixel_data[9][148] = 0;
        pixel_data[9][149] = 0;
        pixel_data[9][150] = 0;
        pixel_data[9][151] = 0;
        pixel_data[9][152] = 0;
        pixel_data[9][153] = 0;
        pixel_data[9][154] = 0;
        pixel_data[9][155] = 0;
        pixel_data[9][156] = 0;
        pixel_data[9][157] = 0;
        pixel_data[9][158] = 0;
        pixel_data[9][159] = 0;
        pixel_data[9][160] = 0;
        pixel_data[9][161] = 0;
        pixel_data[9][162] = 0;
        pixel_data[9][163] = 0;
        pixel_data[9][164] = 0;
        pixel_data[9][165] = 0;
        pixel_data[9][166] = 0;
        pixel_data[9][167] = 0;
        pixel_data[9][168] = 0;
        pixel_data[9][169] = 0;
        pixel_data[9][170] = 0;
        pixel_data[9][171] = 0;
        pixel_data[9][172] = 0;
        pixel_data[9][173] = 0;
        pixel_data[9][174] = 0;
        pixel_data[9][175] = 0;
        pixel_data[9][176] = 0;
        pixel_data[9][177] = 0;
        pixel_data[9][178] = 0;
        pixel_data[9][179] = 0;
        pixel_data[9][180] = 0;
        pixel_data[9][181] = 0;
        pixel_data[9][182] = 0;
        pixel_data[9][183] = 0;
        pixel_data[9][184] = 0;
        pixel_data[9][185] = 0;
        pixel_data[9][186] = 0;
        pixel_data[9][187] = 0;
        pixel_data[9][188] = 0;
        pixel_data[9][189] = 0;
        pixel_data[9][190] = 0;
        pixel_data[9][191] = 0;
        pixel_data[9][192] = 0;
        pixel_data[9][193] = 0;
        pixel_data[9][194] = 0;
        pixel_data[9][195] = 0;
        pixel_data[9][196] = 0;
        pixel_data[9][197] = 0;
        pixel_data[9][198] = 0;
        pixel_data[9][199] = 0; // y=9
        pixel_data[10][0] = 0;
        pixel_data[10][1] = 0;
        pixel_data[10][2] = 0;
        pixel_data[10][3] = 0;
        pixel_data[10][4] = 0;
        pixel_data[10][5] = 0;
        pixel_data[10][6] = 0;
        pixel_data[10][7] = 0;
        pixel_data[10][8] = 0;
        pixel_data[10][9] = 0;
        pixel_data[10][10] = 0;
        pixel_data[10][11] = 0;
        pixel_data[10][12] = 0;
        pixel_data[10][13] = 0;
        pixel_data[10][14] = 0;
        pixel_data[10][15] = 0;
        pixel_data[10][16] = 0;
        pixel_data[10][17] = 0;
        pixel_data[10][18] = 0;
        pixel_data[10][19] = 0;
        pixel_data[10][20] = 0;
        pixel_data[10][21] = 0;
        pixel_data[10][22] = 0;
        pixel_data[10][23] = 0;
        pixel_data[10][24] = 0;
        pixel_data[10][25] = 0;
        pixel_data[10][26] = 0;
        pixel_data[10][27] = 0;
        pixel_data[10][28] = 0;
        pixel_data[10][29] = 0;
        pixel_data[10][30] = 0;
        pixel_data[10][31] = 0;
        pixel_data[10][32] = 0;
        pixel_data[10][33] = 0;
        pixel_data[10][34] = 0;
        pixel_data[10][35] = 0;
        pixel_data[10][36] = 0;
        pixel_data[10][37] = 0;
        pixel_data[10][38] = 0;
        pixel_data[10][39] = 0;
        pixel_data[10][40] = 0;
        pixel_data[10][41] = 0;
        pixel_data[10][42] = 0;
        pixel_data[10][43] = 0;
        pixel_data[10][44] = 0;
        pixel_data[10][45] = 0;
        pixel_data[10][46] = 0;
        pixel_data[10][47] = 0;
        pixel_data[10][48] = 0;
        pixel_data[10][49] = 0;
        pixel_data[10][50] = 0;
        pixel_data[10][51] = 0;
        pixel_data[10][52] = 0;
        pixel_data[10][53] = 0;
        pixel_data[10][54] = 0;
        pixel_data[10][55] = 0;
        pixel_data[10][56] = 0;
        pixel_data[10][57] = 0;
        pixel_data[10][58] = 0;
        pixel_data[10][59] = 0;
        pixel_data[10][60] = 0;
        pixel_data[10][61] = 0;
        pixel_data[10][62] = 0;
        pixel_data[10][63] = 0;
        pixel_data[10][64] = 0;
        pixel_data[10][65] = 0;
        pixel_data[10][66] = 0;
        pixel_data[10][67] = 0;
        pixel_data[10][68] = 0;
        pixel_data[10][69] = 0;
        pixel_data[10][70] = 0;
        pixel_data[10][71] = 0;
        pixel_data[10][72] = 0;
        pixel_data[10][73] = 0;
        pixel_data[10][74] = 0;
        pixel_data[10][75] = 0;
        pixel_data[10][76] = 0;
        pixel_data[10][77] = 0;
        pixel_data[10][78] = 0;
        pixel_data[10][79] = 0;
        pixel_data[10][80] = 0;
        pixel_data[10][81] = 0;
        pixel_data[10][82] = 0;
        pixel_data[10][83] = 0;
        pixel_data[10][84] = 0;
        pixel_data[10][85] = 0;
        pixel_data[10][86] = 0;
        pixel_data[10][87] = 0;
        pixel_data[10][88] = 0;
        pixel_data[10][89] = 0;
        pixel_data[10][90] = 0;
        pixel_data[10][91] = 0;
        pixel_data[10][92] = 0;
        pixel_data[10][93] = 0;
        pixel_data[10][94] = 0;
        pixel_data[10][95] = 0;
        pixel_data[10][96] = 0;
        pixel_data[10][97] = 0;
        pixel_data[10][98] = 0;
        pixel_data[10][99] = 0;
        pixel_data[10][100] = 0;
        pixel_data[10][101] = 0;
        pixel_data[10][102] = 0;
        pixel_data[10][103] = 0;
        pixel_data[10][104] = 0;
        pixel_data[10][105] = 0;
        pixel_data[10][106] = 0;
        pixel_data[10][107] = 0;
        pixel_data[10][108] = 0;
        pixel_data[10][109] = 0;
        pixel_data[10][110] = 0;
        pixel_data[10][111] = 0;
        pixel_data[10][112] = 0;
        pixel_data[10][113] = 0;
        pixel_data[10][114] = 0;
        pixel_data[10][115] = 0;
        pixel_data[10][116] = 0;
        pixel_data[10][117] = 0;
        pixel_data[10][118] = 0;
        pixel_data[10][119] = 0;
        pixel_data[10][120] = 0;
        pixel_data[10][121] = 0;
        pixel_data[10][122] = 0;
        pixel_data[10][123] = 0;
        pixel_data[10][124] = 0;
        pixel_data[10][125] = 0;
        pixel_data[10][126] = 0;
        pixel_data[10][127] = 0;
        pixel_data[10][128] = 0;
        pixel_data[10][129] = 0;
        pixel_data[10][130] = 0;
        pixel_data[10][131] = 0;
        pixel_data[10][132] = 0;
        pixel_data[10][133] = 0;
        pixel_data[10][134] = 0;
        pixel_data[10][135] = 0;
        pixel_data[10][136] = 0;
        pixel_data[10][137] = 0;
        pixel_data[10][138] = 0;
        pixel_data[10][139] = 0;
        pixel_data[10][140] = 0;
        pixel_data[10][141] = 0;
        pixel_data[10][142] = 0;
        pixel_data[10][143] = 0;
        pixel_data[10][144] = 0;
        pixel_data[10][145] = 0;
        pixel_data[10][146] = 0;
        pixel_data[10][147] = 0;
        pixel_data[10][148] = 0;
        pixel_data[10][149] = 0;
        pixel_data[10][150] = 0;
        pixel_data[10][151] = 0;
        pixel_data[10][152] = 0;
        pixel_data[10][153] = 0;
        pixel_data[10][154] = 0;
        pixel_data[10][155] = 0;
        pixel_data[10][156] = 0;
        pixel_data[10][157] = 0;
        pixel_data[10][158] = 0;
        pixel_data[10][159] = 0;
        pixel_data[10][160] = 0;
        pixel_data[10][161] = 0;
        pixel_data[10][162] = 0;
        pixel_data[10][163] = 0;
        pixel_data[10][164] = 0;
        pixel_data[10][165] = 0;
        pixel_data[10][166] = 0;
        pixel_data[10][167] = 0;
        pixel_data[10][168] = 0;
        pixel_data[10][169] = 0;
        pixel_data[10][170] = 0;
        pixel_data[10][171] = 0;
        pixel_data[10][172] = 0;
        pixel_data[10][173] = 0;
        pixel_data[10][174] = 0;
        pixel_data[10][175] = 0;
        pixel_data[10][176] = 0;
        pixel_data[10][177] = 0;
        pixel_data[10][178] = 0;
        pixel_data[10][179] = 0;
        pixel_data[10][180] = 0;
        pixel_data[10][181] = 0;
        pixel_data[10][182] = 0;
        pixel_data[10][183] = 0;
        pixel_data[10][184] = 0;
        pixel_data[10][185] = 0;
        pixel_data[10][186] = 0;
        pixel_data[10][187] = 0;
        pixel_data[10][188] = 0;
        pixel_data[10][189] = 0;
        pixel_data[10][190] = 0;
        pixel_data[10][191] = 0;
        pixel_data[10][192] = 0;
        pixel_data[10][193] = 0;
        pixel_data[10][194] = 0;
        pixel_data[10][195] = 0;
        pixel_data[10][196] = 0;
        pixel_data[10][197] = 0;
        pixel_data[10][198] = 0;
        pixel_data[10][199] = 0; // y=10
        pixel_data[11][0] = 0;
        pixel_data[11][1] = 0;
        pixel_data[11][2] = 0;
        pixel_data[11][3] = 0;
        pixel_data[11][4] = 0;
        pixel_data[11][5] = 0;
        pixel_data[11][6] = 0;
        pixel_data[11][7] = 0;
        pixel_data[11][8] = 0;
        pixel_data[11][9] = 0;
        pixel_data[11][10] = 0;
        pixel_data[11][11] = 0;
        pixel_data[11][12] = 0;
        pixel_data[11][13] = 0;
        pixel_data[11][14] = 0;
        pixel_data[11][15] = 0;
        pixel_data[11][16] = 0;
        pixel_data[11][17] = 0;
        pixel_data[11][18] = 0;
        pixel_data[11][19] = 0;
        pixel_data[11][20] = 0;
        pixel_data[11][21] = 0;
        pixel_data[11][22] = 0;
        pixel_data[11][23] = 0;
        pixel_data[11][24] = 0;
        pixel_data[11][25] = 0;
        pixel_data[11][26] = 0;
        pixel_data[11][27] = 0;
        pixel_data[11][28] = 0;
        pixel_data[11][29] = 0;
        pixel_data[11][30] = 0;
        pixel_data[11][31] = 0;
        pixel_data[11][32] = 0;
        pixel_data[11][33] = 0;
        pixel_data[11][34] = 0;
        pixel_data[11][35] = 0;
        pixel_data[11][36] = 0;
        pixel_data[11][37] = 0;
        pixel_data[11][38] = 0;
        pixel_data[11][39] = 0;
        pixel_data[11][40] = 0;
        pixel_data[11][41] = 0;
        pixel_data[11][42] = 0;
        pixel_data[11][43] = 0;
        pixel_data[11][44] = 0;
        pixel_data[11][45] = 0;
        pixel_data[11][46] = 0;
        pixel_data[11][47] = 0;
        pixel_data[11][48] = 0;
        pixel_data[11][49] = 0;
        pixel_data[11][50] = 0;
        pixel_data[11][51] = 0;
        pixel_data[11][52] = 0;
        pixel_data[11][53] = 0;
        pixel_data[11][54] = 0;
        pixel_data[11][55] = 0;
        pixel_data[11][56] = 0;
        pixel_data[11][57] = 0;
        pixel_data[11][58] = 0;
        pixel_data[11][59] = 0;
        pixel_data[11][60] = 0;
        pixel_data[11][61] = 0;
        pixel_data[11][62] = 0;
        pixel_data[11][63] = 0;
        pixel_data[11][64] = 0;
        pixel_data[11][65] = 0;
        pixel_data[11][66] = 0;
        pixel_data[11][67] = 0;
        pixel_data[11][68] = 0;
        pixel_data[11][69] = 0;
        pixel_data[11][70] = 0;
        pixel_data[11][71] = 0;
        pixel_data[11][72] = 0;
        pixel_data[11][73] = 0;
        pixel_data[11][74] = 0;
        pixel_data[11][75] = 0;
        pixel_data[11][76] = 0;
        pixel_data[11][77] = 0;
        pixel_data[11][78] = 0;
        pixel_data[11][79] = 0;
        pixel_data[11][80] = 0;
        pixel_data[11][81] = 0;
        pixel_data[11][82] = 0;
        pixel_data[11][83] = 0;
        pixel_data[11][84] = 0;
        pixel_data[11][85] = 0;
        pixel_data[11][86] = 0;
        pixel_data[11][87] = 0;
        pixel_data[11][88] = 0;
        pixel_data[11][89] = 0;
        pixel_data[11][90] = 0;
        pixel_data[11][91] = 0;
        pixel_data[11][92] = 0;
        pixel_data[11][93] = 0;
        pixel_data[11][94] = 0;
        pixel_data[11][95] = 0;
        pixel_data[11][96] = 0;
        pixel_data[11][97] = 0;
        pixel_data[11][98] = 0;
        pixel_data[11][99] = 0;
        pixel_data[11][100] = 0;
        pixel_data[11][101] = 0;
        pixel_data[11][102] = 0;
        pixel_data[11][103] = 0;
        pixel_data[11][104] = 0;
        pixel_data[11][105] = 0;
        pixel_data[11][106] = 0;
        pixel_data[11][107] = 0;
        pixel_data[11][108] = 0;
        pixel_data[11][109] = 0;
        pixel_data[11][110] = 0;
        pixel_data[11][111] = 0;
        pixel_data[11][112] = 0;
        pixel_data[11][113] = 0;
        pixel_data[11][114] = 0;
        pixel_data[11][115] = 0;
        pixel_data[11][116] = 0;
        pixel_data[11][117] = 0;
        pixel_data[11][118] = 0;
        pixel_data[11][119] = 0;
        pixel_data[11][120] = 0;
        pixel_data[11][121] = 0;
        pixel_data[11][122] = 0;
        pixel_data[11][123] = 0;
        pixel_data[11][124] = 0;
        pixel_data[11][125] = 0;
        pixel_data[11][126] = 0;
        pixel_data[11][127] = 0;
        pixel_data[11][128] = 0;
        pixel_data[11][129] = 0;
        pixel_data[11][130] = 0;
        pixel_data[11][131] = 0;
        pixel_data[11][132] = 0;
        pixel_data[11][133] = 0;
        pixel_data[11][134] = 0;
        pixel_data[11][135] = 0;
        pixel_data[11][136] = 0;
        pixel_data[11][137] = 0;
        pixel_data[11][138] = 0;
        pixel_data[11][139] = 0;
        pixel_data[11][140] = 0;
        pixel_data[11][141] = 0;
        pixel_data[11][142] = 0;
        pixel_data[11][143] = 0;
        pixel_data[11][144] = 0;
        pixel_data[11][145] = 0;
        pixel_data[11][146] = 0;
        pixel_data[11][147] = 0;
        pixel_data[11][148] = 0;
        pixel_data[11][149] = 0;
        pixel_data[11][150] = 0;
        pixel_data[11][151] = 0;
        pixel_data[11][152] = 0;
        pixel_data[11][153] = 0;
        pixel_data[11][154] = 0;
        pixel_data[11][155] = 0;
        pixel_data[11][156] = 0;
        pixel_data[11][157] = 0;
        pixel_data[11][158] = 0;
        pixel_data[11][159] = 0;
        pixel_data[11][160] = 0;
        pixel_data[11][161] = 0;
        pixel_data[11][162] = 0;
        pixel_data[11][163] = 0;
        pixel_data[11][164] = 0;
        pixel_data[11][165] = 0;
        pixel_data[11][166] = 0;
        pixel_data[11][167] = 0;
        pixel_data[11][168] = 0;
        pixel_data[11][169] = 0;
        pixel_data[11][170] = 0;
        pixel_data[11][171] = 0;
        pixel_data[11][172] = 0;
        pixel_data[11][173] = 0;
        pixel_data[11][174] = 0;
        pixel_data[11][175] = 0;
        pixel_data[11][176] = 0;
        pixel_data[11][177] = 0;
        pixel_data[11][178] = 0;
        pixel_data[11][179] = 0;
        pixel_data[11][180] = 0;
        pixel_data[11][181] = 0;
        pixel_data[11][182] = 0;
        pixel_data[11][183] = 0;
        pixel_data[11][184] = 0;
        pixel_data[11][185] = 0;
        pixel_data[11][186] = 0;
        pixel_data[11][187] = 0;
        pixel_data[11][188] = 0;
        pixel_data[11][189] = 0;
        pixel_data[11][190] = 0;
        pixel_data[11][191] = 0;
        pixel_data[11][192] = 0;
        pixel_data[11][193] = 0;
        pixel_data[11][194] = 0;
        pixel_data[11][195] = 0;
        pixel_data[11][196] = 0;
        pixel_data[11][197] = 0;
        pixel_data[11][198] = 0;
        pixel_data[11][199] = 0; // y=11
        pixel_data[12][0] = 0;
        pixel_data[12][1] = 0;
        pixel_data[12][2] = 0;
        pixel_data[12][3] = 0;
        pixel_data[12][4] = 0;
        pixel_data[12][5] = 0;
        pixel_data[12][6] = 0;
        pixel_data[12][7] = 0;
        pixel_data[12][8] = 0;
        pixel_data[12][9] = 0;
        pixel_data[12][10] = 0;
        pixel_data[12][11] = 0;
        pixel_data[12][12] = 0;
        pixel_data[12][13] = 0;
        pixel_data[12][14] = 0;
        pixel_data[12][15] = 0;
        pixel_data[12][16] = 0;
        pixel_data[12][17] = 0;
        pixel_data[12][18] = 0;
        pixel_data[12][19] = 0;
        pixel_data[12][20] = 0;
        pixel_data[12][21] = 0;
        pixel_data[12][22] = 0;
        pixel_data[12][23] = 0;
        pixel_data[12][24] = 0;
        pixel_data[12][25] = 0;
        pixel_data[12][26] = 0;
        pixel_data[12][27] = 0;
        pixel_data[12][28] = 0;
        pixel_data[12][29] = 0;
        pixel_data[12][30] = 0;
        pixel_data[12][31] = 0;
        pixel_data[12][32] = 0;
        pixel_data[12][33] = 0;
        pixel_data[12][34] = 0;
        pixel_data[12][35] = 0;
        pixel_data[12][36] = 0;
        pixel_data[12][37] = 0;
        pixel_data[12][38] = 0;
        pixel_data[12][39] = 0;
        pixel_data[12][40] = 0;
        pixel_data[12][41] = 0;
        pixel_data[12][42] = 0;
        pixel_data[12][43] = 0;
        pixel_data[12][44] = 0;
        pixel_data[12][45] = 0;
        pixel_data[12][46] = 0;
        pixel_data[12][47] = 0;
        pixel_data[12][48] = 0;
        pixel_data[12][49] = 0;
        pixel_data[12][50] = 0;
        pixel_data[12][51] = 0;
        pixel_data[12][52] = 0;
        pixel_data[12][53] = 0;
        pixel_data[12][54] = 0;
        pixel_data[12][55] = 0;
        pixel_data[12][56] = 0;
        pixel_data[12][57] = 0;
        pixel_data[12][58] = 0;
        pixel_data[12][59] = 0;
        pixel_data[12][60] = 0;
        pixel_data[12][61] = 0;
        pixel_data[12][62] = 0;
        pixel_data[12][63] = 0;
        pixel_data[12][64] = 0;
        pixel_data[12][65] = 0;
        pixel_data[12][66] = 0;
        pixel_data[12][67] = 0;
        pixel_data[12][68] = 0;
        pixel_data[12][69] = 0;
        pixel_data[12][70] = 0;
        pixel_data[12][71] = 0;
        pixel_data[12][72] = 0;
        pixel_data[12][73] = 0;
        pixel_data[12][74] = 0;
        pixel_data[12][75] = 0;
        pixel_data[12][76] = 0;
        pixel_data[12][77] = 0;
        pixel_data[12][78] = 0;
        pixel_data[12][79] = 0;
        pixel_data[12][80] = 0;
        pixel_data[12][81] = 0;
        pixel_data[12][82] = 0;
        pixel_data[12][83] = 0;
        pixel_data[12][84] = 0;
        pixel_data[12][85] = 0;
        pixel_data[12][86] = 0;
        pixel_data[12][87] = 0;
        pixel_data[12][88] = 0;
        pixel_data[12][89] = 0;
        pixel_data[12][90] = 0;
        pixel_data[12][91] = 0;
        pixel_data[12][92] = 0;
        pixel_data[12][93] = 0;
        pixel_data[12][94] = 0;
        pixel_data[12][95] = 0;
        pixel_data[12][96] = 0;
        pixel_data[12][97] = 0;
        pixel_data[12][98] = 0;
        pixel_data[12][99] = 0;
        pixel_data[12][100] = 0;
        pixel_data[12][101] = 0;
        pixel_data[12][102] = 0;
        pixel_data[12][103] = 0;
        pixel_data[12][104] = 0;
        pixel_data[12][105] = 0;
        pixel_data[12][106] = 0;
        pixel_data[12][107] = 0;
        pixel_data[12][108] = 0;
        pixel_data[12][109] = 0;
        pixel_data[12][110] = 0;
        pixel_data[12][111] = 0;
        pixel_data[12][112] = 0;
        pixel_data[12][113] = 0;
        pixel_data[12][114] = 0;
        pixel_data[12][115] = 0;
        pixel_data[12][116] = 0;
        pixel_data[12][117] = 0;
        pixel_data[12][118] = 0;
        pixel_data[12][119] = 0;
        pixel_data[12][120] = 0;
        pixel_data[12][121] = 0;
        pixel_data[12][122] = 0;
        pixel_data[12][123] = 0;
        pixel_data[12][124] = 0;
        pixel_data[12][125] = 0;
        pixel_data[12][126] = 0;
        pixel_data[12][127] = 0;
        pixel_data[12][128] = 0;
        pixel_data[12][129] = 0;
        pixel_data[12][130] = 0;
        pixel_data[12][131] = 0;
        pixel_data[12][132] = 0;
        pixel_data[12][133] = 0;
        pixel_data[12][134] = 0;
        pixel_data[12][135] = 0;
        pixel_data[12][136] = 0;
        pixel_data[12][137] = 0;
        pixel_data[12][138] = 0;
        pixel_data[12][139] = 0;
        pixel_data[12][140] = 0;
        pixel_data[12][141] = 0;
        pixel_data[12][142] = 0;
        pixel_data[12][143] = 0;
        pixel_data[12][144] = 0;
        pixel_data[12][145] = 0;
        pixel_data[12][146] = 0;
        pixel_data[12][147] = 0;
        pixel_data[12][148] = 0;
        pixel_data[12][149] = 0;
        pixel_data[12][150] = 0;
        pixel_data[12][151] = 0;
        pixel_data[12][152] = 0;
        pixel_data[12][153] = 0;
        pixel_data[12][154] = 0;
        pixel_data[12][155] = 0;
        pixel_data[12][156] = 0;
        pixel_data[12][157] = 0;
        pixel_data[12][158] = 0;
        pixel_data[12][159] = 0;
        pixel_data[12][160] = 0;
        pixel_data[12][161] = 0;
        pixel_data[12][162] = 0;
        pixel_data[12][163] = 0;
        pixel_data[12][164] = 0;
        pixel_data[12][165] = 0;
        pixel_data[12][166] = 0;
        pixel_data[12][167] = 0;
        pixel_data[12][168] = 0;
        pixel_data[12][169] = 0;
        pixel_data[12][170] = 0;
        pixel_data[12][171] = 0;
        pixel_data[12][172] = 0;
        pixel_data[12][173] = 0;
        pixel_data[12][174] = 0;
        pixel_data[12][175] = 0;
        pixel_data[12][176] = 0;
        pixel_data[12][177] = 0;
        pixel_data[12][178] = 0;
        pixel_data[12][179] = 0;
        pixel_data[12][180] = 0;
        pixel_data[12][181] = 0;
        pixel_data[12][182] = 0;
        pixel_data[12][183] = 0;
        pixel_data[12][184] = 0;
        pixel_data[12][185] = 0;
        pixel_data[12][186] = 0;
        pixel_data[12][187] = 0;
        pixel_data[12][188] = 0;
        pixel_data[12][189] = 0;
        pixel_data[12][190] = 0;
        pixel_data[12][191] = 0;
        pixel_data[12][192] = 0;
        pixel_data[12][193] = 0;
        pixel_data[12][194] = 0;
        pixel_data[12][195] = 0;
        pixel_data[12][196] = 0;
        pixel_data[12][197] = 0;
        pixel_data[12][198] = 0;
        pixel_data[12][199] = 0; // y=12
        pixel_data[13][0] = 0;
        pixel_data[13][1] = 0;
        pixel_data[13][2] = 0;
        pixel_data[13][3] = 0;
        pixel_data[13][4] = 0;
        pixel_data[13][5] = 0;
        pixel_data[13][6] = 0;
        pixel_data[13][7] = 0;
        pixel_data[13][8] = 0;
        pixel_data[13][9] = 0;
        pixel_data[13][10] = 0;
        pixel_data[13][11] = 0;
        pixel_data[13][12] = 0;
        pixel_data[13][13] = 0;
        pixel_data[13][14] = 0;
        pixel_data[13][15] = 0;
        pixel_data[13][16] = 0;
        pixel_data[13][17] = 0;
        pixel_data[13][18] = 0;
        pixel_data[13][19] = 0;
        pixel_data[13][20] = 0;
        pixel_data[13][21] = 0;
        pixel_data[13][22] = 0;
        pixel_data[13][23] = 0;
        pixel_data[13][24] = 0;
        pixel_data[13][25] = 0;
        pixel_data[13][26] = 0;
        pixel_data[13][27] = 0;
        pixel_data[13][28] = 0;
        pixel_data[13][29] = 0;
        pixel_data[13][30] = 0;
        pixel_data[13][31] = 0;
        pixel_data[13][32] = 0;
        pixel_data[13][33] = 0;
        pixel_data[13][34] = 0;
        pixel_data[13][35] = 0;
        pixel_data[13][36] = 0;
        pixel_data[13][37] = 0;
        pixel_data[13][38] = 0;
        pixel_data[13][39] = 0;
        pixel_data[13][40] = 0;
        pixel_data[13][41] = 0;
        pixel_data[13][42] = 0;
        pixel_data[13][43] = 0;
        pixel_data[13][44] = 0;
        pixel_data[13][45] = 0;
        pixel_data[13][46] = 0;
        pixel_data[13][47] = 0;
        pixel_data[13][48] = 0;
        pixel_data[13][49] = 0;
        pixel_data[13][50] = 0;
        pixel_data[13][51] = 0;
        pixel_data[13][52] = 0;
        pixel_data[13][53] = 0;
        pixel_data[13][54] = 0;
        pixel_data[13][55] = 0;
        pixel_data[13][56] = 0;
        pixel_data[13][57] = 0;
        pixel_data[13][58] = 0;
        pixel_data[13][59] = 0;
        pixel_data[13][60] = 0;
        pixel_data[13][61] = 0;
        pixel_data[13][62] = 0;
        pixel_data[13][63] = 0;
        pixel_data[13][64] = 0;
        pixel_data[13][65] = 0;
        pixel_data[13][66] = 0;
        pixel_data[13][67] = 0;
        pixel_data[13][68] = 0;
        pixel_data[13][69] = 0;
        pixel_data[13][70] = 0;
        pixel_data[13][71] = 0;
        pixel_data[13][72] = 0;
        pixel_data[13][73] = 0;
        pixel_data[13][74] = 0;
        pixel_data[13][75] = 0;
        pixel_data[13][76] = 0;
        pixel_data[13][77] = 0;
        pixel_data[13][78] = 0;
        pixel_data[13][79] = 0;
        pixel_data[13][80] = 0;
        pixel_data[13][81] = 0;
        pixel_data[13][82] = 0;
        pixel_data[13][83] = 0;
        pixel_data[13][84] = 0;
        pixel_data[13][85] = 0;
        pixel_data[13][86] = 0;
        pixel_data[13][87] = 0;
        pixel_data[13][88] = 0;
        pixel_data[13][89] = 0;
        pixel_data[13][90] = 0;
        pixel_data[13][91] = 0;
        pixel_data[13][92] = 0;
        pixel_data[13][93] = 0;
        pixel_data[13][94] = 0;
        pixel_data[13][95] = 0;
        pixel_data[13][96] = 0;
        pixel_data[13][97] = 0;
        pixel_data[13][98] = 0;
        pixel_data[13][99] = 0;
        pixel_data[13][100] = 0;
        pixel_data[13][101] = 0;
        pixel_data[13][102] = 0;
        pixel_data[13][103] = 0;
        pixel_data[13][104] = 0;
        pixel_data[13][105] = 0;
        pixel_data[13][106] = 0;
        pixel_data[13][107] = 0;
        pixel_data[13][108] = 0;
        pixel_data[13][109] = 0;
        pixel_data[13][110] = 0;
        pixel_data[13][111] = 0;
        pixel_data[13][112] = 0;
        pixel_data[13][113] = 0;
        pixel_data[13][114] = 0;
        pixel_data[13][115] = 0;
        pixel_data[13][116] = 0;
        pixel_data[13][117] = 0;
        pixel_data[13][118] = 0;
        pixel_data[13][119] = 0;
        pixel_data[13][120] = 0;
        pixel_data[13][121] = 0;
        pixel_data[13][122] = 0;
        pixel_data[13][123] = 0;
        pixel_data[13][124] = 0;
        pixel_data[13][125] = 0;
        pixel_data[13][126] = 0;
        pixel_data[13][127] = 0;
        pixel_data[13][128] = 0;
        pixel_data[13][129] = 0;
        pixel_data[13][130] = 0;
        pixel_data[13][131] = 0;
        pixel_data[13][132] = 0;
        pixel_data[13][133] = 0;
        pixel_data[13][134] = 0;
        pixel_data[13][135] = 0;
        pixel_data[13][136] = 0;
        pixel_data[13][137] = 0;
        pixel_data[13][138] = 0;
        pixel_data[13][139] = 0;
        pixel_data[13][140] = 0;
        pixel_data[13][141] = 0;
        pixel_data[13][142] = 0;
        pixel_data[13][143] = 0;
        pixel_data[13][144] = 0;
        pixel_data[13][145] = 0;
        pixel_data[13][146] = 0;
        pixel_data[13][147] = 0;
        pixel_data[13][148] = 0;
        pixel_data[13][149] = 0;
        pixel_data[13][150] = 0;
        pixel_data[13][151] = 0;
        pixel_data[13][152] = 0;
        pixel_data[13][153] = 0;
        pixel_data[13][154] = 0;
        pixel_data[13][155] = 0;
        pixel_data[13][156] = 0;
        pixel_data[13][157] = 0;
        pixel_data[13][158] = 0;
        pixel_data[13][159] = 0;
        pixel_data[13][160] = 0;
        pixel_data[13][161] = 0;
        pixel_data[13][162] = 0;
        pixel_data[13][163] = 0;
        pixel_data[13][164] = 0;
        pixel_data[13][165] = 0;
        pixel_data[13][166] = 0;
        pixel_data[13][167] = 0;
        pixel_data[13][168] = 0;
        pixel_data[13][169] = 0;
        pixel_data[13][170] = 0;
        pixel_data[13][171] = 0;
        pixel_data[13][172] = 0;
        pixel_data[13][173] = 0;
        pixel_data[13][174] = 0;
        pixel_data[13][175] = 0;
        pixel_data[13][176] = 0;
        pixel_data[13][177] = 0;
        pixel_data[13][178] = 0;
        pixel_data[13][179] = 0;
        pixel_data[13][180] = 0;
        pixel_data[13][181] = 0;
        pixel_data[13][182] = 0;
        pixel_data[13][183] = 0;
        pixel_data[13][184] = 0;
        pixel_data[13][185] = 0;
        pixel_data[13][186] = 0;
        pixel_data[13][187] = 0;
        pixel_data[13][188] = 0;
        pixel_data[13][189] = 0;
        pixel_data[13][190] = 0;
        pixel_data[13][191] = 0;
        pixel_data[13][192] = 0;
        pixel_data[13][193] = 0;
        pixel_data[13][194] = 0;
        pixel_data[13][195] = 0;
        pixel_data[13][196] = 0;
        pixel_data[13][197] = 0;
        pixel_data[13][198] = 0;
        pixel_data[13][199] = 0; // y=13
        pixel_data[14][0] = 0;
        pixel_data[14][1] = 0;
        pixel_data[14][2] = 0;
        pixel_data[14][3] = 0;
        pixel_data[14][4] = 0;
        pixel_data[14][5] = 0;
        pixel_data[14][6] = 0;
        pixel_data[14][7] = 0;
        pixel_data[14][8] = 0;
        pixel_data[14][9] = 0;
        pixel_data[14][10] = 0;
        pixel_data[14][11] = 0;
        pixel_data[14][12] = 0;
        pixel_data[14][13] = 0;
        pixel_data[14][14] = 0;
        pixel_data[14][15] = 0;
        pixel_data[14][16] = 0;
        pixel_data[14][17] = 0;
        pixel_data[14][18] = 0;
        pixel_data[14][19] = 0;
        pixel_data[14][20] = 0;
        pixel_data[14][21] = 0;
        pixel_data[14][22] = 0;
        pixel_data[14][23] = 0;
        pixel_data[14][24] = 0;
        pixel_data[14][25] = 0;
        pixel_data[14][26] = 0;
        pixel_data[14][27] = 0;
        pixel_data[14][28] = 0;
        pixel_data[14][29] = 0;
        pixel_data[14][30] = 0;
        pixel_data[14][31] = 0;
        pixel_data[14][32] = 0;
        pixel_data[14][33] = 0;
        pixel_data[14][34] = 0;
        pixel_data[14][35] = 0;
        pixel_data[14][36] = 0;
        pixel_data[14][37] = 0;
        pixel_data[14][38] = 0;
        pixel_data[14][39] = 0;
        pixel_data[14][40] = 0;
        pixel_data[14][41] = 0;
        pixel_data[14][42] = 0;
        pixel_data[14][43] = 0;
        pixel_data[14][44] = 0;
        pixel_data[14][45] = 0;
        pixel_data[14][46] = 0;
        pixel_data[14][47] = 0;
        pixel_data[14][48] = 0;
        pixel_data[14][49] = 0;
        pixel_data[14][50] = 0;
        pixel_data[14][51] = 0;
        pixel_data[14][52] = 0;
        pixel_data[14][53] = 0;
        pixel_data[14][54] = 0;
        pixel_data[14][55] = 0;
        pixel_data[14][56] = 0;
        pixel_data[14][57] = 0;
        pixel_data[14][58] = 0;
        pixel_data[14][59] = 0;
        pixel_data[14][60] = 0;
        pixel_data[14][61] = 0;
        pixel_data[14][62] = 0;
        pixel_data[14][63] = 0;
        pixel_data[14][64] = 0;
        pixel_data[14][65] = 0;
        pixel_data[14][66] = 0;
        pixel_data[14][67] = 0;
        pixel_data[14][68] = 0;
        pixel_data[14][69] = 0;
        pixel_data[14][70] = 0;
        pixel_data[14][71] = 0;
        pixel_data[14][72] = 0;
        pixel_data[14][73] = 0;
        pixel_data[14][74] = 0;
        pixel_data[14][75] = 0;
        pixel_data[14][76] = 0;
        pixel_data[14][77] = 0;
        pixel_data[14][78] = 0;
        pixel_data[14][79] = 0;
        pixel_data[14][80] = 0;
        pixel_data[14][81] = 0;
        pixel_data[14][82] = 0;
        pixel_data[14][83] = 0;
        pixel_data[14][84] = 0;
        pixel_data[14][85] = 0;
        pixel_data[14][86] = 0;
        pixel_data[14][87] = 0;
        pixel_data[14][88] = 0;
        pixel_data[14][89] = 0;
        pixel_data[14][90] = 0;
        pixel_data[14][91] = 0;
        pixel_data[14][92] = 0;
        pixel_data[14][93] = 0;
        pixel_data[14][94] = 0;
        pixel_data[14][95] = 0;
        pixel_data[14][96] = 0;
        pixel_data[14][97] = 0;
        pixel_data[14][98] = 0;
        pixel_data[14][99] = 0;
        pixel_data[14][100] = 0;
        pixel_data[14][101] = 0;
        pixel_data[14][102] = 0;
        pixel_data[14][103] = 0;
        pixel_data[14][104] = 0;
        pixel_data[14][105] = 0;
        pixel_data[14][106] = 0;
        pixel_data[14][107] = 0;
        pixel_data[14][108] = 0;
        pixel_data[14][109] = 0;
        pixel_data[14][110] = 0;
        pixel_data[14][111] = 0;
        pixel_data[14][112] = 0;
        pixel_data[14][113] = 0;
        pixel_data[14][114] = 0;
        pixel_data[14][115] = 0;
        pixel_data[14][116] = 0;
        pixel_data[14][117] = 0;
        pixel_data[14][118] = 0;
        pixel_data[14][119] = 0;
        pixel_data[14][120] = 0;
        pixel_data[14][121] = 0;
        pixel_data[14][122] = 0;
        pixel_data[14][123] = 0;
        pixel_data[14][124] = 0;
        pixel_data[14][125] = 0;
        pixel_data[14][126] = 0;
        pixel_data[14][127] = 0;
        pixel_data[14][128] = 0;
        pixel_data[14][129] = 0;
        pixel_data[14][130] = 0;
        pixel_data[14][131] = 0;
        pixel_data[14][132] = 0;
        pixel_data[14][133] = 0;
        pixel_data[14][134] = 0;
        pixel_data[14][135] = 0;
        pixel_data[14][136] = 0;
        pixel_data[14][137] = 0;
        pixel_data[14][138] = 0;
        pixel_data[14][139] = 0;
        pixel_data[14][140] = 0;
        pixel_data[14][141] = 0;
        pixel_data[14][142] = 0;
        pixel_data[14][143] = 0;
        pixel_data[14][144] = 0;
        pixel_data[14][145] = 0;
        pixel_data[14][146] = 0;
        pixel_data[14][147] = 0;
        pixel_data[14][148] = 0;
        pixel_data[14][149] = 0;
        pixel_data[14][150] = 0;
        pixel_data[14][151] = 0;
        pixel_data[14][152] = 0;
        pixel_data[14][153] = 0;
        pixel_data[14][154] = 0;
        pixel_data[14][155] = 0;
        pixel_data[14][156] = 0;
        pixel_data[14][157] = 0;
        pixel_data[14][158] = 0;
        pixel_data[14][159] = 0;
        pixel_data[14][160] = 0;
        pixel_data[14][161] = 0;
        pixel_data[14][162] = 0;
        pixel_data[14][163] = 0;
        pixel_data[14][164] = 0;
        pixel_data[14][165] = 0;
        pixel_data[14][166] = 0;
        pixel_data[14][167] = 0;
        pixel_data[14][168] = 0;
        pixel_data[14][169] = 0;
        pixel_data[14][170] = 0;
        pixel_data[14][171] = 0;
        pixel_data[14][172] = 0;
        pixel_data[14][173] = 0;
        pixel_data[14][174] = 0;
        pixel_data[14][175] = 0;
        pixel_data[14][176] = 0;
        pixel_data[14][177] = 0;
        pixel_data[14][178] = 0;
        pixel_data[14][179] = 0;
        pixel_data[14][180] = 0;
        pixel_data[14][181] = 0;
        pixel_data[14][182] = 0;
        pixel_data[14][183] = 0;
        pixel_data[14][184] = 0;
        pixel_data[14][185] = 0;
        pixel_data[14][186] = 0;
        pixel_data[14][187] = 0;
        pixel_data[14][188] = 0;
        pixel_data[14][189] = 0;
        pixel_data[14][190] = 0;
        pixel_data[14][191] = 0;
        pixel_data[14][192] = 0;
        pixel_data[14][193] = 0;
        pixel_data[14][194] = 0;
        pixel_data[14][195] = 0;
        pixel_data[14][196] = 0;
        pixel_data[14][197] = 0;
        pixel_data[14][198] = 0;
        pixel_data[14][199] = 0; // y=14
        pixel_data[15][0] = 0;
        pixel_data[15][1] = 0;
        pixel_data[15][2] = 0;
        pixel_data[15][3] = 0;
        pixel_data[15][4] = 0;
        pixel_data[15][5] = 0;
        pixel_data[15][6] = 0;
        pixel_data[15][7] = 0;
        pixel_data[15][8] = 0;
        pixel_data[15][9] = 0;
        pixel_data[15][10] = 0;
        pixel_data[15][11] = 0;
        pixel_data[15][12] = 0;
        pixel_data[15][13] = 0;
        pixel_data[15][14] = 0;
        pixel_data[15][15] = 0;
        pixel_data[15][16] = 0;
        pixel_data[15][17] = 0;
        pixel_data[15][18] = 0;
        pixel_data[15][19] = 0;
        pixel_data[15][20] = 0;
        pixel_data[15][21] = 0;
        pixel_data[15][22] = 0;
        pixel_data[15][23] = 0;
        pixel_data[15][24] = 0;
        pixel_data[15][25] = 0;
        pixel_data[15][26] = 0;
        pixel_data[15][27] = 0;
        pixel_data[15][28] = 0;
        pixel_data[15][29] = 0;
        pixel_data[15][30] = 0;
        pixel_data[15][31] = 0;
        pixel_data[15][32] = 0;
        pixel_data[15][33] = 0;
        pixel_data[15][34] = 0;
        pixel_data[15][35] = 0;
        pixel_data[15][36] = 0;
        pixel_data[15][37] = 0;
        pixel_data[15][38] = 0;
        pixel_data[15][39] = 0;
        pixel_data[15][40] = 0;
        pixel_data[15][41] = 0;
        pixel_data[15][42] = 0;
        pixel_data[15][43] = 0;
        pixel_data[15][44] = 0;
        pixel_data[15][45] = 0;
        pixel_data[15][46] = 0;
        pixel_data[15][47] = 0;
        pixel_data[15][48] = 0;
        pixel_data[15][49] = 0;
        pixel_data[15][50] = 0;
        pixel_data[15][51] = 0;
        pixel_data[15][52] = 0;
        pixel_data[15][53] = 0;
        pixel_data[15][54] = 0;
        pixel_data[15][55] = 0;
        pixel_data[15][56] = 0;
        pixel_data[15][57] = 0;
        pixel_data[15][58] = 0;
        pixel_data[15][59] = 0;
        pixel_data[15][60] = 0;
        pixel_data[15][61] = 0;
        pixel_data[15][62] = 0;
        pixel_data[15][63] = 0;
        pixel_data[15][64] = 0;
        pixel_data[15][65] = 0;
        pixel_data[15][66] = 0;
        pixel_data[15][67] = 0;
        pixel_data[15][68] = 0;
        pixel_data[15][69] = 0;
        pixel_data[15][70] = 0;
        pixel_data[15][71] = 0;
        pixel_data[15][72] = 0;
        pixel_data[15][73] = 0;
        pixel_data[15][74] = 0;
        pixel_data[15][75] = 0;
        pixel_data[15][76] = 0;
        pixel_data[15][77] = 0;
        pixel_data[15][78] = 0;
        pixel_data[15][79] = 0;
        pixel_data[15][80] = 0;
        pixel_data[15][81] = 0;
        pixel_data[15][82] = 0;
        pixel_data[15][83] = 0;
        pixel_data[15][84] = 0;
        pixel_data[15][85] = 0;
        pixel_data[15][86] = 0;
        pixel_data[15][87] = 0;
        pixel_data[15][88] = 0;
        pixel_data[15][89] = 0;
        pixel_data[15][90] = 0;
        pixel_data[15][91] = 0;
        pixel_data[15][92] = 0;
        pixel_data[15][93] = 0;
        pixel_data[15][94] = 0;
        pixel_data[15][95] = 0;
        pixel_data[15][96] = 0;
        pixel_data[15][97] = 0;
        pixel_data[15][98] = 0;
        pixel_data[15][99] = 0;
        pixel_data[15][100] = 0;
        pixel_data[15][101] = 0;
        pixel_data[15][102] = 0;
        pixel_data[15][103] = 0;
        pixel_data[15][104] = 0;
        pixel_data[15][105] = 0;
        pixel_data[15][106] = 0;
        pixel_data[15][107] = 0;
        pixel_data[15][108] = 0;
        pixel_data[15][109] = 0;
        pixel_data[15][110] = 0;
        pixel_data[15][111] = 0;
        pixel_data[15][112] = 0;
        pixel_data[15][113] = 0;
        pixel_data[15][114] = 0;
        pixel_data[15][115] = 0;
        pixel_data[15][116] = 0;
        pixel_data[15][117] = 0;
        pixel_data[15][118] = 0;
        pixel_data[15][119] = 0;
        pixel_data[15][120] = 0;
        pixel_data[15][121] = 0;
        pixel_data[15][122] = 0;
        pixel_data[15][123] = 0;
        pixel_data[15][124] = 0;
        pixel_data[15][125] = 0;
        pixel_data[15][126] = 0;
        pixel_data[15][127] = 0;
        pixel_data[15][128] = 0;
        pixel_data[15][129] = 0;
        pixel_data[15][130] = 0;
        pixel_data[15][131] = 0;
        pixel_data[15][132] = 0;
        pixel_data[15][133] = 0;
        pixel_data[15][134] = 0;
        pixel_data[15][135] = 0;
        pixel_data[15][136] = 0;
        pixel_data[15][137] = 0;
        pixel_data[15][138] = 0;
        pixel_data[15][139] = 0;
        pixel_data[15][140] = 0;
        pixel_data[15][141] = 0;
        pixel_data[15][142] = 0;
        pixel_data[15][143] = 0;
        pixel_data[15][144] = 0;
        pixel_data[15][145] = 0;
        pixel_data[15][146] = 0;
        pixel_data[15][147] = 0;
        pixel_data[15][148] = 0;
        pixel_data[15][149] = 0;
        pixel_data[15][150] = 0;
        pixel_data[15][151] = 0;
        pixel_data[15][152] = 0;
        pixel_data[15][153] = 0;
        pixel_data[15][154] = 0;
        pixel_data[15][155] = 0;
        pixel_data[15][156] = 0;
        pixel_data[15][157] = 0;
        pixel_data[15][158] = 0;
        pixel_data[15][159] = 0;
        pixel_data[15][160] = 0;
        pixel_data[15][161] = 0;
        pixel_data[15][162] = 0;
        pixel_data[15][163] = 0;
        pixel_data[15][164] = 0;
        pixel_data[15][165] = 0;
        pixel_data[15][166] = 0;
        pixel_data[15][167] = 0;
        pixel_data[15][168] = 0;
        pixel_data[15][169] = 0;
        pixel_data[15][170] = 0;
        pixel_data[15][171] = 0;
        pixel_data[15][172] = 0;
        pixel_data[15][173] = 0;
        pixel_data[15][174] = 0;
        pixel_data[15][175] = 0;
        pixel_data[15][176] = 0;
        pixel_data[15][177] = 0;
        pixel_data[15][178] = 0;
        pixel_data[15][179] = 0;
        pixel_data[15][180] = 0;
        pixel_data[15][181] = 0;
        pixel_data[15][182] = 0;
        pixel_data[15][183] = 0;
        pixel_data[15][184] = 0;
        pixel_data[15][185] = 0;
        pixel_data[15][186] = 0;
        pixel_data[15][187] = 0;
        pixel_data[15][188] = 0;
        pixel_data[15][189] = 0;
        pixel_data[15][190] = 0;
        pixel_data[15][191] = 0;
        pixel_data[15][192] = 0;
        pixel_data[15][193] = 0;
        pixel_data[15][194] = 0;
        pixel_data[15][195] = 0;
        pixel_data[15][196] = 0;
        pixel_data[15][197] = 0;
        pixel_data[15][198] = 0;
        pixel_data[15][199] = 0; // y=15
        pixel_data[16][0] = 0;
        pixel_data[16][1] = 0;
        pixel_data[16][2] = 0;
        pixel_data[16][3] = 0;
        pixel_data[16][4] = 0;
        pixel_data[16][5] = 0;
        pixel_data[16][6] = 0;
        pixel_data[16][7] = 0;
        pixel_data[16][8] = 0;
        pixel_data[16][9] = 0;
        pixel_data[16][10] = 0;
        pixel_data[16][11] = 0;
        pixel_data[16][12] = 0;
        pixel_data[16][13] = 0;
        pixel_data[16][14] = 0;
        pixel_data[16][15] = 0;
        pixel_data[16][16] = 0;
        pixel_data[16][17] = 0;
        pixel_data[16][18] = 0;
        pixel_data[16][19] = 0;
        pixel_data[16][20] = 0;
        pixel_data[16][21] = 0;
        pixel_data[16][22] = 0;
        pixel_data[16][23] = 0;
        pixel_data[16][24] = 0;
        pixel_data[16][25] = 0;
        pixel_data[16][26] = 0;
        pixel_data[16][27] = 0;
        pixel_data[16][28] = 0;
        pixel_data[16][29] = 0;
        pixel_data[16][30] = 0;
        pixel_data[16][31] = 0;
        pixel_data[16][32] = 0;
        pixel_data[16][33] = 0;
        pixel_data[16][34] = 0;
        pixel_data[16][35] = 0;
        pixel_data[16][36] = 0;
        pixel_data[16][37] = 0;
        pixel_data[16][38] = 0;
        pixel_data[16][39] = 0;
        pixel_data[16][40] = 0;
        pixel_data[16][41] = 0;
        pixel_data[16][42] = 0;
        pixel_data[16][43] = 0;
        pixel_data[16][44] = 0;
        pixel_data[16][45] = 0;
        pixel_data[16][46] = 0;
        pixel_data[16][47] = 0;
        pixel_data[16][48] = 0;
        pixel_data[16][49] = 0;
        pixel_data[16][50] = 0;
        pixel_data[16][51] = 0;
        pixel_data[16][52] = 0;
        pixel_data[16][53] = 0;
        pixel_data[16][54] = 0;
        pixel_data[16][55] = 0;
        pixel_data[16][56] = 0;
        pixel_data[16][57] = 0;
        pixel_data[16][58] = 0;
        pixel_data[16][59] = 0;
        pixel_data[16][60] = 0;
        pixel_data[16][61] = 0;
        pixel_data[16][62] = 0;
        pixel_data[16][63] = 0;
        pixel_data[16][64] = 0;
        pixel_data[16][65] = 0;
        pixel_data[16][66] = 0;
        pixel_data[16][67] = 0;
        pixel_data[16][68] = 0;
        pixel_data[16][69] = 0;
        pixel_data[16][70] = 0;
        pixel_data[16][71] = 0;
        pixel_data[16][72] = 0;
        pixel_data[16][73] = 0;
        pixel_data[16][74] = 0;
        pixel_data[16][75] = 0;
        pixel_data[16][76] = 0;
        pixel_data[16][77] = 0;
        pixel_data[16][78] = 0;
        pixel_data[16][79] = 0;
        pixel_data[16][80] = 0;
        pixel_data[16][81] = 0;
        pixel_data[16][82] = 0;
        pixel_data[16][83] = 0;
        pixel_data[16][84] = 0;
        pixel_data[16][85] = 0;
        pixel_data[16][86] = 0;
        pixel_data[16][87] = 0;
        pixel_data[16][88] = 0;
        pixel_data[16][89] = 0;
        pixel_data[16][90] = 0;
        pixel_data[16][91] = 0;
        pixel_data[16][92] = 0;
        pixel_data[16][93] = 0;
        pixel_data[16][94] = 0;
        pixel_data[16][95] = 0;
        pixel_data[16][96] = 0;
        pixel_data[16][97] = 0;
        pixel_data[16][98] = 0;
        pixel_data[16][99] = 0;
        pixel_data[16][100] = 0;
        pixel_data[16][101] = 0;
        pixel_data[16][102] = 0;
        pixel_data[16][103] = 0;
        pixel_data[16][104] = 0;
        pixel_data[16][105] = 0;
        pixel_data[16][106] = 0;
        pixel_data[16][107] = 0;
        pixel_data[16][108] = 0;
        pixel_data[16][109] = 0;
        pixel_data[16][110] = 0;
        pixel_data[16][111] = 0;
        pixel_data[16][112] = 0;
        pixel_data[16][113] = 0;
        pixel_data[16][114] = 0;
        pixel_data[16][115] = 0;
        pixel_data[16][116] = 0;
        pixel_data[16][117] = 0;
        pixel_data[16][118] = 0;
        pixel_data[16][119] = 0;
        pixel_data[16][120] = 0;
        pixel_data[16][121] = 0;
        pixel_data[16][122] = 0;
        pixel_data[16][123] = 0;
        pixel_data[16][124] = 0;
        pixel_data[16][125] = 0;
        pixel_data[16][126] = 0;
        pixel_data[16][127] = 0;
        pixel_data[16][128] = 0;
        pixel_data[16][129] = 0;
        pixel_data[16][130] = 0;
        pixel_data[16][131] = 0;
        pixel_data[16][132] = 0;
        pixel_data[16][133] = 0;
        pixel_data[16][134] = 0;
        pixel_data[16][135] = 0;
        pixel_data[16][136] = 0;
        pixel_data[16][137] = 0;
        pixel_data[16][138] = 0;
        pixel_data[16][139] = 0;
        pixel_data[16][140] = 0;
        pixel_data[16][141] = 0;
        pixel_data[16][142] = 0;
        pixel_data[16][143] = 0;
        pixel_data[16][144] = 0;
        pixel_data[16][145] = 0;
        pixel_data[16][146] = 0;
        pixel_data[16][147] = 0;
        pixel_data[16][148] = 0;
        pixel_data[16][149] = 0;
        pixel_data[16][150] = 0;
        pixel_data[16][151] = 0;
        pixel_data[16][152] = 0;
        pixel_data[16][153] = 0;
        pixel_data[16][154] = 0;
        pixel_data[16][155] = 0;
        pixel_data[16][156] = 0;
        pixel_data[16][157] = 0;
        pixel_data[16][158] = 0;
        pixel_data[16][159] = 0;
        pixel_data[16][160] = 0;
        pixel_data[16][161] = 0;
        pixel_data[16][162] = 0;
        pixel_data[16][163] = 0;
        pixel_data[16][164] = 0;
        pixel_data[16][165] = 0;
        pixel_data[16][166] = 0;
        pixel_data[16][167] = 0;
        pixel_data[16][168] = 0;
        pixel_data[16][169] = 0;
        pixel_data[16][170] = 0;
        pixel_data[16][171] = 0;
        pixel_data[16][172] = 0;
        pixel_data[16][173] = 0;
        pixel_data[16][174] = 0;
        pixel_data[16][175] = 0;
        pixel_data[16][176] = 0;
        pixel_data[16][177] = 0;
        pixel_data[16][178] = 0;
        pixel_data[16][179] = 0;
        pixel_data[16][180] = 0;
        pixel_data[16][181] = 0;
        pixel_data[16][182] = 0;
        pixel_data[16][183] = 0;
        pixel_data[16][184] = 0;
        pixel_data[16][185] = 0;
        pixel_data[16][186] = 0;
        pixel_data[16][187] = 0;
        pixel_data[16][188] = 0;
        pixel_data[16][189] = 0;
        pixel_data[16][190] = 0;
        pixel_data[16][191] = 0;
        pixel_data[16][192] = 0;
        pixel_data[16][193] = 0;
        pixel_data[16][194] = 0;
        pixel_data[16][195] = 0;
        pixel_data[16][196] = 0;
        pixel_data[16][197] = 0;
        pixel_data[16][198] = 0;
        pixel_data[16][199] = 0; // y=16
        pixel_data[17][0] = 0;
        pixel_data[17][1] = 0;
        pixel_data[17][2] = 0;
        pixel_data[17][3] = 0;
        pixel_data[17][4] = 0;
        pixel_data[17][5] = 0;
        pixel_data[17][6] = 0;
        pixel_data[17][7] = 0;
        pixel_data[17][8] = 0;
        pixel_data[17][9] = 0;
        pixel_data[17][10] = 0;
        pixel_data[17][11] = 0;
        pixel_data[17][12] = 0;
        pixel_data[17][13] = 0;
        pixel_data[17][14] = 0;
        pixel_data[17][15] = 0;
        pixel_data[17][16] = 0;
        pixel_data[17][17] = 0;
        pixel_data[17][18] = 0;
        pixel_data[17][19] = 0;
        pixel_data[17][20] = 0;
        pixel_data[17][21] = 0;
        pixel_data[17][22] = 0;
        pixel_data[17][23] = 0;
        pixel_data[17][24] = 0;
        pixel_data[17][25] = 0;
        pixel_data[17][26] = 0;
        pixel_data[17][27] = 0;
        pixel_data[17][28] = 0;
        pixel_data[17][29] = 0;
        pixel_data[17][30] = 0;
        pixel_data[17][31] = 0;
        pixel_data[17][32] = 0;
        pixel_data[17][33] = 0;
        pixel_data[17][34] = 0;
        pixel_data[17][35] = 0;
        pixel_data[17][36] = 0;
        pixel_data[17][37] = 0;
        pixel_data[17][38] = 0;
        pixel_data[17][39] = 0;
        pixel_data[17][40] = 0;
        pixel_data[17][41] = 0;
        pixel_data[17][42] = 0;
        pixel_data[17][43] = 0;
        pixel_data[17][44] = 0;
        pixel_data[17][45] = 0;
        pixel_data[17][46] = 0;
        pixel_data[17][47] = 0;
        pixel_data[17][48] = 0;
        pixel_data[17][49] = 0;
        pixel_data[17][50] = 0;
        pixel_data[17][51] = 0;
        pixel_data[17][52] = 0;
        pixel_data[17][53] = 0;
        pixel_data[17][54] = 0;
        pixel_data[17][55] = 0;
        pixel_data[17][56] = 0;
        pixel_data[17][57] = 0;
        pixel_data[17][58] = 0;
        pixel_data[17][59] = 0;
        pixel_data[17][60] = 0;
        pixel_data[17][61] = 0;
        pixel_data[17][62] = 0;
        pixel_data[17][63] = 0;
        pixel_data[17][64] = 0;
        pixel_data[17][65] = 0;
        pixel_data[17][66] = 0;
        pixel_data[17][67] = 0;
        pixel_data[17][68] = 0;
        pixel_data[17][69] = 0;
        pixel_data[17][70] = 0;
        pixel_data[17][71] = 0;
        pixel_data[17][72] = 0;
        pixel_data[17][73] = 0;
        pixel_data[17][74] = 0;
        pixel_data[17][75] = 0;
        pixel_data[17][76] = 0;
        pixel_data[17][77] = 0;
        pixel_data[17][78] = 0;
        pixel_data[17][79] = 0;
        pixel_data[17][80] = 0;
        pixel_data[17][81] = 0;
        pixel_data[17][82] = 0;
        pixel_data[17][83] = 0;
        pixel_data[17][84] = 0;
        pixel_data[17][85] = 0;
        pixel_data[17][86] = 0;
        pixel_data[17][87] = 0;
        pixel_data[17][88] = 0;
        pixel_data[17][89] = 0;
        pixel_data[17][90] = 0;
        pixel_data[17][91] = 0;
        pixel_data[17][92] = 0;
        pixel_data[17][93] = 0;
        pixel_data[17][94] = 0;
        pixel_data[17][95] = 0;
        pixel_data[17][96] = 0;
        pixel_data[17][97] = 0;
        pixel_data[17][98] = 0;
        pixel_data[17][99] = 0;
        pixel_data[17][100] = 0;
        pixel_data[17][101] = 0;
        pixel_data[17][102] = 0;
        pixel_data[17][103] = 0;
        pixel_data[17][104] = 0;
        pixel_data[17][105] = 0;
        pixel_data[17][106] = 0;
        pixel_data[17][107] = 0;
        pixel_data[17][108] = 0;
        pixel_data[17][109] = 0;
        pixel_data[17][110] = 0;
        pixel_data[17][111] = 0;
        pixel_data[17][112] = 0;
        pixel_data[17][113] = 0;
        pixel_data[17][114] = 0;
        pixel_data[17][115] = 0;
        pixel_data[17][116] = 0;
        pixel_data[17][117] = 0;
        pixel_data[17][118] = 0;
        pixel_data[17][119] = 0;
        pixel_data[17][120] = 0;
        pixel_data[17][121] = 0;
        pixel_data[17][122] = 0;
        pixel_data[17][123] = 0;
        pixel_data[17][124] = 0;
        pixel_data[17][125] = 0;
        pixel_data[17][126] = 0;
        pixel_data[17][127] = 0;
        pixel_data[17][128] = 0;
        pixel_data[17][129] = 0;
        pixel_data[17][130] = 0;
        pixel_data[17][131] = 0;
        pixel_data[17][132] = 0;
        pixel_data[17][133] = 0;
        pixel_data[17][134] = 0;
        pixel_data[17][135] = 0;
        pixel_data[17][136] = 0;
        pixel_data[17][137] = 0;
        pixel_data[17][138] = 0;
        pixel_data[17][139] = 0;
        pixel_data[17][140] = 0;
        pixel_data[17][141] = 0;
        pixel_data[17][142] = 0;
        pixel_data[17][143] = 0;
        pixel_data[17][144] = 0;
        pixel_data[17][145] = 0;
        pixel_data[17][146] = 0;
        pixel_data[17][147] = 0;
        pixel_data[17][148] = 0;
        pixel_data[17][149] = 0;
        pixel_data[17][150] = 0;
        pixel_data[17][151] = 0;
        pixel_data[17][152] = 0;
        pixel_data[17][153] = 0;
        pixel_data[17][154] = 0;
        pixel_data[17][155] = 0;
        pixel_data[17][156] = 0;
        pixel_data[17][157] = 0;
        pixel_data[17][158] = 0;
        pixel_data[17][159] = 0;
        pixel_data[17][160] = 0;
        pixel_data[17][161] = 0;
        pixel_data[17][162] = 0;
        pixel_data[17][163] = 0;
        pixel_data[17][164] = 0;
        pixel_data[17][165] = 0;
        pixel_data[17][166] = 0;
        pixel_data[17][167] = 0;
        pixel_data[17][168] = 0;
        pixel_data[17][169] = 0;
        pixel_data[17][170] = 0;
        pixel_data[17][171] = 0;
        pixel_data[17][172] = 0;
        pixel_data[17][173] = 0;
        pixel_data[17][174] = 0;
        pixel_data[17][175] = 0;
        pixel_data[17][176] = 0;
        pixel_data[17][177] = 0;
        pixel_data[17][178] = 0;
        pixel_data[17][179] = 0;
        pixel_data[17][180] = 0;
        pixel_data[17][181] = 0;
        pixel_data[17][182] = 0;
        pixel_data[17][183] = 0;
        pixel_data[17][184] = 0;
        pixel_data[17][185] = 0;
        pixel_data[17][186] = 0;
        pixel_data[17][187] = 0;
        pixel_data[17][188] = 0;
        pixel_data[17][189] = 0;
        pixel_data[17][190] = 0;
        pixel_data[17][191] = 0;
        pixel_data[17][192] = 0;
        pixel_data[17][193] = 0;
        pixel_data[17][194] = 0;
        pixel_data[17][195] = 0;
        pixel_data[17][196] = 0;
        pixel_data[17][197] = 0;
        pixel_data[17][198] = 0;
        pixel_data[17][199] = 0; // y=17
        pixel_data[18][0] = 0;
        pixel_data[18][1] = 0;
        pixel_data[18][2] = 0;
        pixel_data[18][3] = 0;
        pixel_data[18][4] = 0;
        pixel_data[18][5] = 0;
        pixel_data[18][6] = 0;
        pixel_data[18][7] = 0;
        pixel_data[18][8] = 0;
        pixel_data[18][9] = 0;
        pixel_data[18][10] = 0;
        pixel_data[18][11] = 0;
        pixel_data[18][12] = 0;
        pixel_data[18][13] = 0;
        pixel_data[18][14] = 0;
        pixel_data[18][15] = 0;
        pixel_data[18][16] = 0;
        pixel_data[18][17] = 0;
        pixel_data[18][18] = 0;
        pixel_data[18][19] = 0;
        pixel_data[18][20] = 0;
        pixel_data[18][21] = 0;
        pixel_data[18][22] = 0;
        pixel_data[18][23] = 0;
        pixel_data[18][24] = 0;
        pixel_data[18][25] = 0;
        pixel_data[18][26] = 0;
        pixel_data[18][27] = 0;
        pixel_data[18][28] = 0;
        pixel_data[18][29] = 0;
        pixel_data[18][30] = 0;
        pixel_data[18][31] = 0;
        pixel_data[18][32] = 0;
        pixel_data[18][33] = 0;
        pixel_data[18][34] = 0;
        pixel_data[18][35] = 0;
        pixel_data[18][36] = 0;
        pixel_data[18][37] = 0;
        pixel_data[18][38] = 0;
        pixel_data[18][39] = 0;
        pixel_data[18][40] = 0;
        pixel_data[18][41] = 0;
        pixel_data[18][42] = 0;
        pixel_data[18][43] = 0;
        pixel_data[18][44] = 0;
        pixel_data[18][45] = 0;
        pixel_data[18][46] = 0;
        pixel_data[18][47] = 0;
        pixel_data[18][48] = 0;
        pixel_data[18][49] = 0;
        pixel_data[18][50] = 0;
        pixel_data[18][51] = 0;
        pixel_data[18][52] = 0;
        pixel_data[18][53] = 0;
        pixel_data[18][54] = 0;
        pixel_data[18][55] = 0;
        pixel_data[18][56] = 0;
        pixel_data[18][57] = 0;
        pixel_data[18][58] = 0;
        pixel_data[18][59] = 0;
        pixel_data[18][60] = 0;
        pixel_data[18][61] = 0;
        pixel_data[18][62] = 0;
        pixel_data[18][63] = 0;
        pixel_data[18][64] = 0;
        pixel_data[18][65] = 0;
        pixel_data[18][66] = 0;
        pixel_data[18][67] = 0;
        pixel_data[18][68] = 0;
        pixel_data[18][69] = 0;
        pixel_data[18][70] = 0;
        pixel_data[18][71] = 0;
        pixel_data[18][72] = 0;
        pixel_data[18][73] = 0;
        pixel_data[18][74] = 0;
        pixel_data[18][75] = 0;
        pixel_data[18][76] = 0;
        pixel_data[18][77] = 0;
        pixel_data[18][78] = 0;
        pixel_data[18][79] = 0;
        pixel_data[18][80] = 0;
        pixel_data[18][81] = 0;
        pixel_data[18][82] = 0;
        pixel_data[18][83] = 0;
        pixel_data[18][84] = 0;
        pixel_data[18][85] = 0;
        pixel_data[18][86] = 0;
        pixel_data[18][87] = 0;
        pixel_data[18][88] = 0;
        pixel_data[18][89] = 0;
        pixel_data[18][90] = 0;
        pixel_data[18][91] = 0;
        pixel_data[18][92] = 0;
        pixel_data[18][93] = 0;
        pixel_data[18][94] = 0;
        pixel_data[18][95] = 0;
        pixel_data[18][96] = 0;
        pixel_data[18][97] = 0;
        pixel_data[18][98] = 0;
        pixel_data[18][99] = 0;
        pixel_data[18][100] = 0;
        pixel_data[18][101] = 0;
        pixel_data[18][102] = 0;
        pixel_data[18][103] = 0;
        pixel_data[18][104] = 0;
        pixel_data[18][105] = 0;
        pixel_data[18][106] = 0;
        pixel_data[18][107] = 0;
        pixel_data[18][108] = 0;
        pixel_data[18][109] = 0;
        pixel_data[18][110] = 0;
        pixel_data[18][111] = 0;
        pixel_data[18][112] = 0;
        pixel_data[18][113] = 0;
        pixel_data[18][114] = 0;
        pixel_data[18][115] = 0;
        pixel_data[18][116] = 0;
        pixel_data[18][117] = 0;
        pixel_data[18][118] = 0;
        pixel_data[18][119] = 0;
        pixel_data[18][120] = 0;
        pixel_data[18][121] = 0;
        pixel_data[18][122] = 0;
        pixel_data[18][123] = 0;
        pixel_data[18][124] = 0;
        pixel_data[18][125] = 0;
        pixel_data[18][126] = 0;
        pixel_data[18][127] = 0;
        pixel_data[18][128] = 0;
        pixel_data[18][129] = 0;
        pixel_data[18][130] = 0;
        pixel_data[18][131] = 0;
        pixel_data[18][132] = 0;
        pixel_data[18][133] = 0;
        pixel_data[18][134] = 0;
        pixel_data[18][135] = 0;
        pixel_data[18][136] = 0;
        pixel_data[18][137] = 0;
        pixel_data[18][138] = 0;
        pixel_data[18][139] = 0;
        pixel_data[18][140] = 0;
        pixel_data[18][141] = 0;
        pixel_data[18][142] = 0;
        pixel_data[18][143] = 0;
        pixel_data[18][144] = 0;
        pixel_data[18][145] = 0;
        pixel_data[18][146] = 0;
        pixel_data[18][147] = 0;
        pixel_data[18][148] = 0;
        pixel_data[18][149] = 0;
        pixel_data[18][150] = 0;
        pixel_data[18][151] = 0;
        pixel_data[18][152] = 0;
        pixel_data[18][153] = 0;
        pixel_data[18][154] = 0;
        pixel_data[18][155] = 0;
        pixel_data[18][156] = 0;
        pixel_data[18][157] = 0;
        pixel_data[18][158] = 0;
        pixel_data[18][159] = 0;
        pixel_data[18][160] = 0;
        pixel_data[18][161] = 0;
        pixel_data[18][162] = 0;
        pixel_data[18][163] = 0;
        pixel_data[18][164] = 0;
        pixel_data[18][165] = 0;
        pixel_data[18][166] = 0;
        pixel_data[18][167] = 0;
        pixel_data[18][168] = 0;
        pixel_data[18][169] = 0;
        pixel_data[18][170] = 0;
        pixel_data[18][171] = 0;
        pixel_data[18][172] = 0;
        pixel_data[18][173] = 0;
        pixel_data[18][174] = 0;
        pixel_data[18][175] = 0;
        pixel_data[18][176] = 0;
        pixel_data[18][177] = 0;
        pixel_data[18][178] = 0;
        pixel_data[18][179] = 0;
        pixel_data[18][180] = 0;
        pixel_data[18][181] = 0;
        pixel_data[18][182] = 0;
        pixel_data[18][183] = 0;
        pixel_data[18][184] = 0;
        pixel_data[18][185] = 0;
        pixel_data[18][186] = 0;
        pixel_data[18][187] = 0;
        pixel_data[18][188] = 0;
        pixel_data[18][189] = 0;
        pixel_data[18][190] = 0;
        pixel_data[18][191] = 0;
        pixel_data[18][192] = 0;
        pixel_data[18][193] = 0;
        pixel_data[18][194] = 0;
        pixel_data[18][195] = 0;
        pixel_data[18][196] = 0;
        pixel_data[18][197] = 0;
        pixel_data[18][198] = 0;
        pixel_data[18][199] = 0; // y=18
        pixel_data[19][0] = 0;
        pixel_data[19][1] = 0;
        pixel_data[19][2] = 0;
        pixel_data[19][3] = 0;
        pixel_data[19][4] = 0;
        pixel_data[19][5] = 0;
        pixel_data[19][6] = 0;
        pixel_data[19][7] = 0;
        pixel_data[19][8] = 0;
        pixel_data[19][9] = 0;
        pixel_data[19][10] = 0;
        pixel_data[19][11] = 0;
        pixel_data[19][12] = 0;
        pixel_data[19][13] = 0;
        pixel_data[19][14] = 0;
        pixel_data[19][15] = 0;
        pixel_data[19][16] = 0;
        pixel_data[19][17] = 0;
        pixel_data[19][18] = 0;
        pixel_data[19][19] = 0;
        pixel_data[19][20] = 0;
        pixel_data[19][21] = 0;
        pixel_data[19][22] = 0;
        pixel_data[19][23] = 0;
        pixel_data[19][24] = 0;
        pixel_data[19][25] = 0;
        pixel_data[19][26] = 0;
        pixel_data[19][27] = 0;
        pixel_data[19][28] = 0;
        pixel_data[19][29] = 0;
        pixel_data[19][30] = 0;
        pixel_data[19][31] = 0;
        pixel_data[19][32] = 0;
        pixel_data[19][33] = 0;
        pixel_data[19][34] = 0;
        pixel_data[19][35] = 0;
        pixel_data[19][36] = 0;
        pixel_data[19][37] = 0;
        pixel_data[19][38] = 0;
        pixel_data[19][39] = 0;
        pixel_data[19][40] = 0;
        pixel_data[19][41] = 0;
        pixel_data[19][42] = 0;
        pixel_data[19][43] = 0;
        pixel_data[19][44] = 0;
        pixel_data[19][45] = 0;
        pixel_data[19][46] = 0;
        pixel_data[19][47] = 0;
        pixel_data[19][48] = 0;
        pixel_data[19][49] = 0;
        pixel_data[19][50] = 0;
        pixel_data[19][51] = 0;
        pixel_data[19][52] = 0;
        pixel_data[19][53] = 0;
        pixel_data[19][54] = 0;
        pixel_data[19][55] = 0;
        pixel_data[19][56] = 0;
        pixel_data[19][57] = 0;
        pixel_data[19][58] = 0;
        pixel_data[19][59] = 0;
        pixel_data[19][60] = 0;
        pixel_data[19][61] = 0;
        pixel_data[19][62] = 0;
        pixel_data[19][63] = 0;
        pixel_data[19][64] = 0;
        pixel_data[19][65] = 0;
        pixel_data[19][66] = 0;
        pixel_data[19][67] = 0;
        pixel_data[19][68] = 0;
        pixel_data[19][69] = 0;
        pixel_data[19][70] = 0;
        pixel_data[19][71] = 0;
        pixel_data[19][72] = 0;
        pixel_data[19][73] = 0;
        pixel_data[19][74] = 0;
        pixel_data[19][75] = 0;
        pixel_data[19][76] = 0;
        pixel_data[19][77] = 0;
        pixel_data[19][78] = 0;
        pixel_data[19][79] = 0;
        pixel_data[19][80] = 0;
        pixel_data[19][81] = 0;
        pixel_data[19][82] = 0;
        pixel_data[19][83] = 0;
        pixel_data[19][84] = 0;
        pixel_data[19][85] = 0;
        pixel_data[19][86] = 0;
        pixel_data[19][87] = 0;
        pixel_data[19][88] = 0;
        pixel_data[19][89] = 0;
        pixel_data[19][90] = 0;
        pixel_data[19][91] = 0;
        pixel_data[19][92] = 0;
        pixel_data[19][93] = 0;
        pixel_data[19][94] = 0;
        pixel_data[19][95] = 0;
        pixel_data[19][96] = 0;
        pixel_data[19][97] = 0;
        pixel_data[19][98] = 0;
        pixel_data[19][99] = 0;
        pixel_data[19][100] = 0;
        pixel_data[19][101] = 0;
        pixel_data[19][102] = 0;
        pixel_data[19][103] = 0;
        pixel_data[19][104] = 0;
        pixel_data[19][105] = 0;
        pixel_data[19][106] = 0;
        pixel_data[19][107] = 0;
        pixel_data[19][108] = 0;
        pixel_data[19][109] = 0;
        pixel_data[19][110] = 0;
        pixel_data[19][111] = 0;
        pixel_data[19][112] = 0;
        pixel_data[19][113] = 0;
        pixel_data[19][114] = 0;
        pixel_data[19][115] = 0;
        pixel_data[19][116] = 0;
        pixel_data[19][117] = 0;
        pixel_data[19][118] = 0;
        pixel_data[19][119] = 0;
        pixel_data[19][120] = 0;
        pixel_data[19][121] = 0;
        pixel_data[19][122] = 0;
        pixel_data[19][123] = 0;
        pixel_data[19][124] = 0;
        pixel_data[19][125] = 0;
        pixel_data[19][126] = 0;
        pixel_data[19][127] = 0;
        pixel_data[19][128] = 0;
        pixel_data[19][129] = 0;
        pixel_data[19][130] = 0;
        pixel_data[19][131] = 0;
        pixel_data[19][132] = 0;
        pixel_data[19][133] = 0;
        pixel_data[19][134] = 0;
        pixel_data[19][135] = 0;
        pixel_data[19][136] = 0;
        pixel_data[19][137] = 0;
        pixel_data[19][138] = 0;
        pixel_data[19][139] = 0;
        pixel_data[19][140] = 0;
        pixel_data[19][141] = 0;
        pixel_data[19][142] = 0;
        pixel_data[19][143] = 0;
        pixel_data[19][144] = 0;
        pixel_data[19][145] = 0;
        pixel_data[19][146] = 0;
        pixel_data[19][147] = 0;
        pixel_data[19][148] = 0;
        pixel_data[19][149] = 0;
        pixel_data[19][150] = 0;
        pixel_data[19][151] = 0;
        pixel_data[19][152] = 0;
        pixel_data[19][153] = 0;
        pixel_data[19][154] = 0;
        pixel_data[19][155] = 0;
        pixel_data[19][156] = 0;
        pixel_data[19][157] = 0;
        pixel_data[19][158] = 0;
        pixel_data[19][159] = 0;
        pixel_data[19][160] = 0;
        pixel_data[19][161] = 0;
        pixel_data[19][162] = 0;
        pixel_data[19][163] = 0;
        pixel_data[19][164] = 0;
        pixel_data[19][165] = 0;
        pixel_data[19][166] = 0;
        pixel_data[19][167] = 0;
        pixel_data[19][168] = 0;
        pixel_data[19][169] = 0;
        pixel_data[19][170] = 0;
        pixel_data[19][171] = 0;
        pixel_data[19][172] = 0;
        pixel_data[19][173] = 0;
        pixel_data[19][174] = 0;
        pixel_data[19][175] = 0;
        pixel_data[19][176] = 0;
        pixel_data[19][177] = 0;
        pixel_data[19][178] = 0;
        pixel_data[19][179] = 0;
        pixel_data[19][180] = 0;
        pixel_data[19][181] = 0;
        pixel_data[19][182] = 0;
        pixel_data[19][183] = 0;
        pixel_data[19][184] = 0;
        pixel_data[19][185] = 0;
        pixel_data[19][186] = 0;
        pixel_data[19][187] = 0;
        pixel_data[19][188] = 0;
        pixel_data[19][189] = 0;
        pixel_data[19][190] = 0;
        pixel_data[19][191] = 0;
        pixel_data[19][192] = 0;
        pixel_data[19][193] = 0;
        pixel_data[19][194] = 0;
        pixel_data[19][195] = 0;
        pixel_data[19][196] = 0;
        pixel_data[19][197] = 0;
        pixel_data[19][198] = 0;
        pixel_data[19][199] = 0; // y=19
        pixel_data[20][0] = 0;
        pixel_data[20][1] = 0;
        pixel_data[20][2] = 0;
        pixel_data[20][3] = 0;
        pixel_data[20][4] = 0;
        pixel_data[20][5] = 0;
        pixel_data[20][6] = 0;
        pixel_data[20][7] = 0;
        pixel_data[20][8] = 0;
        pixel_data[20][9] = 0;
        pixel_data[20][10] = 0;
        pixel_data[20][11] = 0;
        pixel_data[20][12] = 0;
        pixel_data[20][13] = 0;
        pixel_data[20][14] = 0;
        pixel_data[20][15] = 0;
        pixel_data[20][16] = 0;
        pixel_data[20][17] = 0;
        pixel_data[20][18] = 0;
        pixel_data[20][19] = 0;
        pixel_data[20][20] = 0;
        pixel_data[20][21] = 0;
        pixel_data[20][22] = 0;
        pixel_data[20][23] = 0;
        pixel_data[20][24] = 0;
        pixel_data[20][25] = 0;
        pixel_data[20][26] = 0;
        pixel_data[20][27] = 0;
        pixel_data[20][28] = 0;
        pixel_data[20][29] = 0;
        pixel_data[20][30] = 0;
        pixel_data[20][31] = 0;
        pixel_data[20][32] = 0;
        pixel_data[20][33] = 0;
        pixel_data[20][34] = 0;
        pixel_data[20][35] = 0;
        pixel_data[20][36] = 0;
        pixel_data[20][37] = 0;
        pixel_data[20][38] = 0;
        pixel_data[20][39] = 0;
        pixel_data[20][40] = 0;
        pixel_data[20][41] = 0;
        pixel_data[20][42] = 0;
        pixel_data[20][43] = 0;
        pixel_data[20][44] = 0;
        pixel_data[20][45] = 0;
        pixel_data[20][46] = 0;
        pixel_data[20][47] = 0;
        pixel_data[20][48] = 0;
        pixel_data[20][49] = 0;
        pixel_data[20][50] = 0;
        pixel_data[20][51] = 0;
        pixel_data[20][52] = 0;
        pixel_data[20][53] = 0;
        pixel_data[20][54] = 0;
        pixel_data[20][55] = 0;
        pixel_data[20][56] = 0;
        pixel_data[20][57] = 0;
        pixel_data[20][58] = 0;
        pixel_data[20][59] = 0;
        pixel_data[20][60] = 0;
        pixel_data[20][61] = 0;
        pixel_data[20][62] = 0;
        pixel_data[20][63] = 0;
        pixel_data[20][64] = 0;
        pixel_data[20][65] = 0;
        pixel_data[20][66] = 0;
        pixel_data[20][67] = 0;
        pixel_data[20][68] = 0;
        pixel_data[20][69] = 0;
        pixel_data[20][70] = 0;
        pixel_data[20][71] = 0;
        pixel_data[20][72] = 0;
        pixel_data[20][73] = 0;
        pixel_data[20][74] = 0;
        pixel_data[20][75] = 0;
        pixel_data[20][76] = 0;
        pixel_data[20][77] = 0;
        pixel_data[20][78] = 0;
        pixel_data[20][79] = 0;
        pixel_data[20][80] = 0;
        pixel_data[20][81] = 0;
        pixel_data[20][82] = 0;
        pixel_data[20][83] = 0;
        pixel_data[20][84] = 0;
        pixel_data[20][85] = 0;
        pixel_data[20][86] = 0;
        pixel_data[20][87] = 0;
        pixel_data[20][88] = 0;
        pixel_data[20][89] = 0;
        pixel_data[20][90] = 0;
        pixel_data[20][91] = 0;
        pixel_data[20][92] = 0;
        pixel_data[20][93] = 0;
        pixel_data[20][94] = 0;
        pixel_data[20][95] = 0;
        pixel_data[20][96] = 0;
        pixel_data[20][97] = 0;
        pixel_data[20][98] = 0;
        pixel_data[20][99] = 0;
        pixel_data[20][100] = 0;
        pixel_data[20][101] = 0;
        pixel_data[20][102] = 0;
        pixel_data[20][103] = 0;
        pixel_data[20][104] = 0;
        pixel_data[20][105] = 0;
        pixel_data[20][106] = 0;
        pixel_data[20][107] = 0;
        pixel_data[20][108] = 0;
        pixel_data[20][109] = 0;
        pixel_data[20][110] = 0;
        pixel_data[20][111] = 0;
        pixel_data[20][112] = 0;
        pixel_data[20][113] = 0;
        pixel_data[20][114] = 0;
        pixel_data[20][115] = 0;
        pixel_data[20][116] = 0;
        pixel_data[20][117] = 0;
        pixel_data[20][118] = 0;
        pixel_data[20][119] = 0;
        pixel_data[20][120] = 0;
        pixel_data[20][121] = 0;
        pixel_data[20][122] = 0;
        pixel_data[20][123] = 0;
        pixel_data[20][124] = 0;
        pixel_data[20][125] = 0;
        pixel_data[20][126] = 0;
        pixel_data[20][127] = 0;
        pixel_data[20][128] = 0;
        pixel_data[20][129] = 0;
        pixel_data[20][130] = 0;
        pixel_data[20][131] = 0;
        pixel_data[20][132] = 0;
        pixel_data[20][133] = 0;
        pixel_data[20][134] = 0;
        pixel_data[20][135] = 0;
        pixel_data[20][136] = 0;
        pixel_data[20][137] = 0;
        pixel_data[20][138] = 0;
        pixel_data[20][139] = 0;
        pixel_data[20][140] = 0;
        pixel_data[20][141] = 0;
        pixel_data[20][142] = 0;
        pixel_data[20][143] = 0;
        pixel_data[20][144] = 0;
        pixel_data[20][145] = 0;
        pixel_data[20][146] = 0;
        pixel_data[20][147] = 0;
        pixel_data[20][148] = 0;
        pixel_data[20][149] = 0;
        pixel_data[20][150] = 0;
        pixel_data[20][151] = 0;
        pixel_data[20][152] = 0;
        pixel_data[20][153] = 0;
        pixel_data[20][154] = 0;
        pixel_data[20][155] = 0;
        pixel_data[20][156] = 0;
        pixel_data[20][157] = 0;
        pixel_data[20][158] = 0;
        pixel_data[20][159] = 0;
        pixel_data[20][160] = 0;
        pixel_data[20][161] = 0;
        pixel_data[20][162] = 0;
        pixel_data[20][163] = 0;
        pixel_data[20][164] = 0;
        pixel_data[20][165] = 0;
        pixel_data[20][166] = 0;
        pixel_data[20][167] = 0;
        pixel_data[20][168] = 0;
        pixel_data[20][169] = 0;
        pixel_data[20][170] = 0;
        pixel_data[20][171] = 0;
        pixel_data[20][172] = 0;
        pixel_data[20][173] = 0;
        pixel_data[20][174] = 0;
        pixel_data[20][175] = 0;
        pixel_data[20][176] = 0;
        pixel_data[20][177] = 0;
        pixel_data[20][178] = 0;
        pixel_data[20][179] = 0;
        pixel_data[20][180] = 0;
        pixel_data[20][181] = 0;
        pixel_data[20][182] = 0;
        pixel_data[20][183] = 0;
        pixel_data[20][184] = 0;
        pixel_data[20][185] = 0;
        pixel_data[20][186] = 0;
        pixel_data[20][187] = 0;
        pixel_data[20][188] = 0;
        pixel_data[20][189] = 0;
        pixel_data[20][190] = 0;
        pixel_data[20][191] = 0;
        pixel_data[20][192] = 0;
        pixel_data[20][193] = 0;
        pixel_data[20][194] = 0;
        pixel_data[20][195] = 0;
        pixel_data[20][196] = 0;
        pixel_data[20][197] = 0;
        pixel_data[20][198] = 0;
        pixel_data[20][199] = 0; // y=20
        pixel_data[21][0] = 0;
        pixel_data[21][1] = 0;
        pixel_data[21][2] = 0;
        pixel_data[21][3] = 0;
        pixel_data[21][4] = 0;
        pixel_data[21][5] = 0;
        pixel_data[21][6] = 0;
        pixel_data[21][7] = 0;
        pixel_data[21][8] = 0;
        pixel_data[21][9] = 0;
        pixel_data[21][10] = 0;
        pixel_data[21][11] = 0;
        pixel_data[21][12] = 0;
        pixel_data[21][13] = 0;
        pixel_data[21][14] = 0;
        pixel_data[21][15] = 0;
        pixel_data[21][16] = 0;
        pixel_data[21][17] = 0;
        pixel_data[21][18] = 0;
        pixel_data[21][19] = 0;
        pixel_data[21][20] = 0;
        pixel_data[21][21] = 0;
        pixel_data[21][22] = 0;
        pixel_data[21][23] = 0;
        pixel_data[21][24] = 0;
        pixel_data[21][25] = 0;
        pixel_data[21][26] = 0;
        pixel_data[21][27] = 0;
        pixel_data[21][28] = 0;
        pixel_data[21][29] = 0;
        pixel_data[21][30] = 0;
        pixel_data[21][31] = 0;
        pixel_data[21][32] = 0;
        pixel_data[21][33] = 0;
        pixel_data[21][34] = 0;
        pixel_data[21][35] = 0;
        pixel_data[21][36] = 0;
        pixel_data[21][37] = 0;
        pixel_data[21][38] = 0;
        pixel_data[21][39] = 0;
        pixel_data[21][40] = 0;
        pixel_data[21][41] = 0;
        pixel_data[21][42] = 0;
        pixel_data[21][43] = 0;
        pixel_data[21][44] = 0;
        pixel_data[21][45] = 0;
        pixel_data[21][46] = 0;
        pixel_data[21][47] = 0;
        pixel_data[21][48] = 0;
        pixel_data[21][49] = 0;
        pixel_data[21][50] = 0;
        pixel_data[21][51] = 0;
        pixel_data[21][52] = 0;
        pixel_data[21][53] = 0;
        pixel_data[21][54] = 0;
        pixel_data[21][55] = 0;
        pixel_data[21][56] = 0;
        pixel_data[21][57] = 0;
        pixel_data[21][58] = 0;
        pixel_data[21][59] = 0;
        pixel_data[21][60] = 0;
        pixel_data[21][61] = 0;
        pixel_data[21][62] = 0;
        pixel_data[21][63] = 0;
        pixel_data[21][64] = 0;
        pixel_data[21][65] = 0;
        pixel_data[21][66] = 0;
        pixel_data[21][67] = 0;
        pixel_data[21][68] = 0;
        pixel_data[21][69] = 0;
        pixel_data[21][70] = 0;
        pixel_data[21][71] = 0;
        pixel_data[21][72] = 0;
        pixel_data[21][73] = 0;
        pixel_data[21][74] = 0;
        pixel_data[21][75] = 0;
        pixel_data[21][76] = 0;
        pixel_data[21][77] = 0;
        pixel_data[21][78] = 0;
        pixel_data[21][79] = 0;
        pixel_data[21][80] = 0;
        pixel_data[21][81] = 0;
        pixel_data[21][82] = 0;
        pixel_data[21][83] = 0;
        pixel_data[21][84] = 0;
        pixel_data[21][85] = 0;
        pixel_data[21][86] = 0;
        pixel_data[21][87] = 0;
        pixel_data[21][88] = 0;
        pixel_data[21][89] = 0;
        pixel_data[21][90] = 0;
        pixel_data[21][91] = 0;
        pixel_data[21][92] = 0;
        pixel_data[21][93] = 0;
        pixel_data[21][94] = 0;
        pixel_data[21][95] = 0;
        pixel_data[21][96] = 0;
        pixel_data[21][97] = 0;
        pixel_data[21][98] = 0;
        pixel_data[21][99] = 0;
        pixel_data[21][100] = 0;
        pixel_data[21][101] = 0;
        pixel_data[21][102] = 0;
        pixel_data[21][103] = 0;
        pixel_data[21][104] = 0;
        pixel_data[21][105] = 0;
        pixel_data[21][106] = 0;
        pixel_data[21][107] = 0;
        pixel_data[21][108] = 0;
        pixel_data[21][109] = 0;
        pixel_data[21][110] = 0;
        pixel_data[21][111] = 0;
        pixel_data[21][112] = 0;
        pixel_data[21][113] = 0;
        pixel_data[21][114] = 0;
        pixel_data[21][115] = 0;
        pixel_data[21][116] = 0;
        pixel_data[21][117] = 0;
        pixel_data[21][118] = 0;
        pixel_data[21][119] = 0;
        pixel_data[21][120] = 0;
        pixel_data[21][121] = 0;
        pixel_data[21][122] = 0;
        pixel_data[21][123] = 0;
        pixel_data[21][124] = 0;
        pixel_data[21][125] = 0;
        pixel_data[21][126] = 0;
        pixel_data[21][127] = 0;
        pixel_data[21][128] = 0;
        pixel_data[21][129] = 0;
        pixel_data[21][130] = 0;
        pixel_data[21][131] = 0;
        pixel_data[21][132] = 0;
        pixel_data[21][133] = 0;
        pixel_data[21][134] = 0;
        pixel_data[21][135] = 0;
        pixel_data[21][136] = 0;
        pixel_data[21][137] = 0;
        pixel_data[21][138] = 0;
        pixel_data[21][139] = 0;
        pixel_data[21][140] = 0;
        pixel_data[21][141] = 0;
        pixel_data[21][142] = 0;
        pixel_data[21][143] = 0;
        pixel_data[21][144] = 0;
        pixel_data[21][145] = 0;
        pixel_data[21][146] = 0;
        pixel_data[21][147] = 0;
        pixel_data[21][148] = 0;
        pixel_data[21][149] = 0;
        pixel_data[21][150] = 0;
        pixel_data[21][151] = 0;
        pixel_data[21][152] = 0;
        pixel_data[21][153] = 0;
        pixel_data[21][154] = 0;
        pixel_data[21][155] = 0;
        pixel_data[21][156] = 0;
        pixel_data[21][157] = 0;
        pixel_data[21][158] = 0;
        pixel_data[21][159] = 0;
        pixel_data[21][160] = 0;
        pixel_data[21][161] = 0;
        pixel_data[21][162] = 0;
        pixel_data[21][163] = 0;
        pixel_data[21][164] = 0;
        pixel_data[21][165] = 0;
        pixel_data[21][166] = 0;
        pixel_data[21][167] = 0;
        pixel_data[21][168] = 0;
        pixel_data[21][169] = 0;
        pixel_data[21][170] = 0;
        pixel_data[21][171] = 0;
        pixel_data[21][172] = 0;
        pixel_data[21][173] = 0;
        pixel_data[21][174] = 0;
        pixel_data[21][175] = 0;
        pixel_data[21][176] = 0;
        pixel_data[21][177] = 0;
        pixel_data[21][178] = 0;
        pixel_data[21][179] = 0;
        pixel_data[21][180] = 0;
        pixel_data[21][181] = 0;
        pixel_data[21][182] = 0;
        pixel_data[21][183] = 0;
        pixel_data[21][184] = 0;
        pixel_data[21][185] = 0;
        pixel_data[21][186] = 0;
        pixel_data[21][187] = 0;
        pixel_data[21][188] = 0;
        pixel_data[21][189] = 0;
        pixel_data[21][190] = 0;
        pixel_data[21][191] = 0;
        pixel_data[21][192] = 0;
        pixel_data[21][193] = 0;
        pixel_data[21][194] = 0;
        pixel_data[21][195] = 0;
        pixel_data[21][196] = 0;
        pixel_data[21][197] = 0;
        pixel_data[21][198] = 0;
        pixel_data[21][199] = 0; // y=21
        pixel_data[22][0] = 0;
        pixel_data[22][1] = 0;
        pixel_data[22][2] = 0;
        pixel_data[22][3] = 0;
        pixel_data[22][4] = 0;
        pixel_data[22][5] = 0;
        pixel_data[22][6] = 0;
        pixel_data[22][7] = 0;
        pixel_data[22][8] = 0;
        pixel_data[22][9] = 0;
        pixel_data[22][10] = 0;
        pixel_data[22][11] = 0;
        pixel_data[22][12] = 0;
        pixel_data[22][13] = 0;
        pixel_data[22][14] = 0;
        pixel_data[22][15] = 0;
        pixel_data[22][16] = 0;
        pixel_data[22][17] = 0;
        pixel_data[22][18] = 0;
        pixel_data[22][19] = 0;
        pixel_data[22][20] = 0;
        pixel_data[22][21] = 0;
        pixel_data[22][22] = 0;
        pixel_data[22][23] = 0;
        pixel_data[22][24] = 0;
        pixel_data[22][25] = 0;
        pixel_data[22][26] = 0;
        pixel_data[22][27] = 0;
        pixel_data[22][28] = 0;
        pixel_data[22][29] = 0;
        pixel_data[22][30] = 0;
        pixel_data[22][31] = 0;
        pixel_data[22][32] = 0;
        pixel_data[22][33] = 0;
        pixel_data[22][34] = 0;
        pixel_data[22][35] = 0;
        pixel_data[22][36] = 0;
        pixel_data[22][37] = 0;
        pixel_data[22][38] = 0;
        pixel_data[22][39] = 0;
        pixel_data[22][40] = 0;
        pixel_data[22][41] = 0;
        pixel_data[22][42] = 0;
        pixel_data[22][43] = 0;
        pixel_data[22][44] = 0;
        pixel_data[22][45] = 0;
        pixel_data[22][46] = 0;
        pixel_data[22][47] = 0;
        pixel_data[22][48] = 0;
        pixel_data[22][49] = 0;
        pixel_data[22][50] = 0;
        pixel_data[22][51] = 0;
        pixel_data[22][52] = 0;
        pixel_data[22][53] = 0;
        pixel_data[22][54] = 0;
        pixel_data[22][55] = 0;
        pixel_data[22][56] = 0;
        pixel_data[22][57] = 0;
        pixel_data[22][58] = 0;
        pixel_data[22][59] = 0;
        pixel_data[22][60] = 0;
        pixel_data[22][61] = 0;
        pixel_data[22][62] = 0;
        pixel_data[22][63] = 0;
        pixel_data[22][64] = 0;
        pixel_data[22][65] = 0;
        pixel_data[22][66] = 0;
        pixel_data[22][67] = 0;
        pixel_data[22][68] = 0;
        pixel_data[22][69] = 0;
        pixel_data[22][70] = 0;
        pixel_data[22][71] = 0;
        pixel_data[22][72] = 0;
        pixel_data[22][73] = 0;
        pixel_data[22][74] = 0;
        pixel_data[22][75] = 0;
        pixel_data[22][76] = 0;
        pixel_data[22][77] = 0;
        pixel_data[22][78] = 0;
        pixel_data[22][79] = 0;
        pixel_data[22][80] = 0;
        pixel_data[22][81] = 0;
        pixel_data[22][82] = 0;
        pixel_data[22][83] = 0;
        pixel_data[22][84] = 0;
        pixel_data[22][85] = 0;
        pixel_data[22][86] = 0;
        pixel_data[22][87] = 0;
        pixel_data[22][88] = 0;
        pixel_data[22][89] = 0;
        pixel_data[22][90] = 0;
        pixel_data[22][91] = 0;
        pixel_data[22][92] = 0;
        pixel_data[22][93] = 0;
        pixel_data[22][94] = 0;
        pixel_data[22][95] = 0;
        pixel_data[22][96] = 0;
        pixel_data[22][97] = 0;
        pixel_data[22][98] = 0;
        pixel_data[22][99] = 0;
        pixel_data[22][100] = 0;
        pixel_data[22][101] = 0;
        pixel_data[22][102] = 0;
        pixel_data[22][103] = 0;
        pixel_data[22][104] = 0;
        pixel_data[22][105] = 0;
        pixel_data[22][106] = 0;
        pixel_data[22][107] = 0;
        pixel_data[22][108] = 0;
        pixel_data[22][109] = 0;
        pixel_data[22][110] = 0;
        pixel_data[22][111] = 0;
        pixel_data[22][112] = 0;
        pixel_data[22][113] = 0;
        pixel_data[22][114] = 0;
        pixel_data[22][115] = 0;
        pixel_data[22][116] = 0;
        pixel_data[22][117] = 0;
        pixel_data[22][118] = 0;
        pixel_data[22][119] = 0;
        pixel_data[22][120] = 0;
        pixel_data[22][121] = 0;
        pixel_data[22][122] = 0;
        pixel_data[22][123] = 0;
        pixel_data[22][124] = 0;
        pixel_data[22][125] = 0;
        pixel_data[22][126] = 0;
        pixel_data[22][127] = 0;
        pixel_data[22][128] = 0;
        pixel_data[22][129] = 0;
        pixel_data[22][130] = 0;
        pixel_data[22][131] = 0;
        pixel_data[22][132] = 0;
        pixel_data[22][133] = 0;
        pixel_data[22][134] = 0;
        pixel_data[22][135] = 0;
        pixel_data[22][136] = 0;
        pixel_data[22][137] = 0;
        pixel_data[22][138] = 0;
        pixel_data[22][139] = 0;
        pixel_data[22][140] = 0;
        pixel_data[22][141] = 0;
        pixel_data[22][142] = 0;
        pixel_data[22][143] = 0;
        pixel_data[22][144] = 0;
        pixel_data[22][145] = 0;
        pixel_data[22][146] = 0;
        pixel_data[22][147] = 0;
        pixel_data[22][148] = 0;
        pixel_data[22][149] = 0;
        pixel_data[22][150] = 0;
        pixel_data[22][151] = 0;
        pixel_data[22][152] = 0;
        pixel_data[22][153] = 0;
        pixel_data[22][154] = 0;
        pixel_data[22][155] = 0;
        pixel_data[22][156] = 0;
        pixel_data[22][157] = 0;
        pixel_data[22][158] = 0;
        pixel_data[22][159] = 0;
        pixel_data[22][160] = 0;
        pixel_data[22][161] = 0;
        pixel_data[22][162] = 0;
        pixel_data[22][163] = 0;
        pixel_data[22][164] = 0;
        pixel_data[22][165] = 0;
        pixel_data[22][166] = 0;
        pixel_data[22][167] = 0;
        pixel_data[22][168] = 0;
        pixel_data[22][169] = 0;
        pixel_data[22][170] = 0;
        pixel_data[22][171] = 0;
        pixel_data[22][172] = 0;
        pixel_data[22][173] = 0;
        pixel_data[22][174] = 0;
        pixel_data[22][175] = 0;
        pixel_data[22][176] = 0;
        pixel_data[22][177] = 0;
        pixel_data[22][178] = 0;
        pixel_data[22][179] = 0;
        pixel_data[22][180] = 0;
        pixel_data[22][181] = 0;
        pixel_data[22][182] = 0;
        pixel_data[22][183] = 0;
        pixel_data[22][184] = 0;
        pixel_data[22][185] = 0;
        pixel_data[22][186] = 0;
        pixel_data[22][187] = 0;
        pixel_data[22][188] = 0;
        pixel_data[22][189] = 0;
        pixel_data[22][190] = 0;
        pixel_data[22][191] = 0;
        pixel_data[22][192] = 0;
        pixel_data[22][193] = 0;
        pixel_data[22][194] = 0;
        pixel_data[22][195] = 0;
        pixel_data[22][196] = 0;
        pixel_data[22][197] = 0;
        pixel_data[22][198] = 0;
        pixel_data[22][199] = 0; // y=22
        pixel_data[23][0] = 0;
        pixel_data[23][1] = 0;
        pixel_data[23][2] = 0;
        pixel_data[23][3] = 0;
        pixel_data[23][4] = 0;
        pixel_data[23][5] = 0;
        pixel_data[23][6] = 0;
        pixel_data[23][7] = 0;
        pixel_data[23][8] = 0;
        pixel_data[23][9] = 0;
        pixel_data[23][10] = 0;
        pixel_data[23][11] = 0;
        pixel_data[23][12] = 0;
        pixel_data[23][13] = 0;
        pixel_data[23][14] = 0;
        pixel_data[23][15] = 0;
        pixel_data[23][16] = 0;
        pixel_data[23][17] = 0;
        pixel_data[23][18] = 0;
        pixel_data[23][19] = 0;
        pixel_data[23][20] = 0;
        pixel_data[23][21] = 0;
        pixel_data[23][22] = 0;
        pixel_data[23][23] = 0;
        pixel_data[23][24] = 0;
        pixel_data[23][25] = 0;
        pixel_data[23][26] = 0;
        pixel_data[23][27] = 0;
        pixel_data[23][28] = 0;
        pixel_data[23][29] = 0;
        pixel_data[23][30] = 0;
        pixel_data[23][31] = 0;
        pixel_data[23][32] = 0;
        pixel_data[23][33] = 0;
        pixel_data[23][34] = 0;
        pixel_data[23][35] = 0;
        pixel_data[23][36] = 0;
        pixel_data[23][37] = 0;
        pixel_data[23][38] = 0;
        pixel_data[23][39] = 0;
        pixel_data[23][40] = 0;
        pixel_data[23][41] = 0;
        pixel_data[23][42] = 0;
        pixel_data[23][43] = 0;
        pixel_data[23][44] = 0;
        pixel_data[23][45] = 0;
        pixel_data[23][46] = 0;
        pixel_data[23][47] = 0;
        pixel_data[23][48] = 0;
        pixel_data[23][49] = 0;
        pixel_data[23][50] = 0;
        pixel_data[23][51] = 0;
        pixel_data[23][52] = 0;
        pixel_data[23][53] = 0;
        pixel_data[23][54] = 0;
        pixel_data[23][55] = 0;
        pixel_data[23][56] = 0;
        pixel_data[23][57] = 0;
        pixel_data[23][58] = 0;
        pixel_data[23][59] = 0;
        pixel_data[23][60] = 0;
        pixel_data[23][61] = 0;
        pixel_data[23][62] = 0;
        pixel_data[23][63] = 0;
        pixel_data[23][64] = 0;
        pixel_data[23][65] = 0;
        pixel_data[23][66] = 0;
        pixel_data[23][67] = 0;
        pixel_data[23][68] = 0;
        pixel_data[23][69] = 0;
        pixel_data[23][70] = 0;
        pixel_data[23][71] = 0;
        pixel_data[23][72] = 0;
        pixel_data[23][73] = 0;
        pixel_data[23][74] = 0;
        pixel_data[23][75] = 0;
        pixel_data[23][76] = 0;
        pixel_data[23][77] = 0;
        pixel_data[23][78] = 0;
        pixel_data[23][79] = 0;
        pixel_data[23][80] = 0;
        pixel_data[23][81] = 0;
        pixel_data[23][82] = 0;
        pixel_data[23][83] = 0;
        pixel_data[23][84] = 0;
        pixel_data[23][85] = 0;
        pixel_data[23][86] = 0;
        pixel_data[23][87] = 0;
        pixel_data[23][88] = 0;
        pixel_data[23][89] = 0;
        pixel_data[23][90] = 0;
        pixel_data[23][91] = 0;
        pixel_data[23][92] = 0;
        pixel_data[23][93] = 0;
        pixel_data[23][94] = 0;
        pixel_data[23][95] = 0;
        pixel_data[23][96] = 0;
        pixel_data[23][97] = 0;
        pixel_data[23][98] = 0;
        pixel_data[23][99] = 0;
        pixel_data[23][100] = 0;
        pixel_data[23][101] = 0;
        pixel_data[23][102] = 0;
        pixel_data[23][103] = 0;
        pixel_data[23][104] = 0;
        pixel_data[23][105] = 0;
        pixel_data[23][106] = 0;
        pixel_data[23][107] = 0;
        pixel_data[23][108] = 0;
        pixel_data[23][109] = 0;
        pixel_data[23][110] = 0;
        pixel_data[23][111] = 0;
        pixel_data[23][112] = 0;
        pixel_data[23][113] = 0;
        pixel_data[23][114] = 0;
        pixel_data[23][115] = 0;
        pixel_data[23][116] = 0;
        pixel_data[23][117] = 0;
        pixel_data[23][118] = 0;
        pixel_data[23][119] = 0;
        pixel_data[23][120] = 0;
        pixel_data[23][121] = 0;
        pixel_data[23][122] = 0;
        pixel_data[23][123] = 0;
        pixel_data[23][124] = 0;
        pixel_data[23][125] = 0;
        pixel_data[23][126] = 0;
        pixel_data[23][127] = 0;
        pixel_data[23][128] = 0;
        pixel_data[23][129] = 0;
        pixel_data[23][130] = 0;
        pixel_data[23][131] = 0;
        pixel_data[23][132] = 0;
        pixel_data[23][133] = 0;
        pixel_data[23][134] = 0;
        pixel_data[23][135] = 0;
        pixel_data[23][136] = 0;
        pixel_data[23][137] = 0;
        pixel_data[23][138] = 0;
        pixel_data[23][139] = 0;
        pixel_data[23][140] = 0;
        pixel_data[23][141] = 0;
        pixel_data[23][142] = 0;
        pixel_data[23][143] = 0;
        pixel_data[23][144] = 0;
        pixel_data[23][145] = 0;
        pixel_data[23][146] = 0;
        pixel_data[23][147] = 0;
        pixel_data[23][148] = 0;
        pixel_data[23][149] = 0;
        pixel_data[23][150] = 0;
        pixel_data[23][151] = 0;
        pixel_data[23][152] = 0;
        pixel_data[23][153] = 0;
        pixel_data[23][154] = 0;
        pixel_data[23][155] = 0;
        pixel_data[23][156] = 0;
        pixel_data[23][157] = 0;
        pixel_data[23][158] = 0;
        pixel_data[23][159] = 0;
        pixel_data[23][160] = 0;
        pixel_data[23][161] = 0;
        pixel_data[23][162] = 0;
        pixel_data[23][163] = 0;
        pixel_data[23][164] = 0;
        pixel_data[23][165] = 0;
        pixel_data[23][166] = 0;
        pixel_data[23][167] = 0;
        pixel_data[23][168] = 0;
        pixel_data[23][169] = 0;
        pixel_data[23][170] = 0;
        pixel_data[23][171] = 0;
        pixel_data[23][172] = 0;
        pixel_data[23][173] = 0;
        pixel_data[23][174] = 0;
        pixel_data[23][175] = 0;
        pixel_data[23][176] = 0;
        pixel_data[23][177] = 0;
        pixel_data[23][178] = 0;
        pixel_data[23][179] = 0;
        pixel_data[23][180] = 0;
        pixel_data[23][181] = 0;
        pixel_data[23][182] = 0;
        pixel_data[23][183] = 0;
        pixel_data[23][184] = 0;
        pixel_data[23][185] = 0;
        pixel_data[23][186] = 0;
        pixel_data[23][187] = 0;
        pixel_data[23][188] = 0;
        pixel_data[23][189] = 0;
        pixel_data[23][190] = 0;
        pixel_data[23][191] = 0;
        pixel_data[23][192] = 0;
        pixel_data[23][193] = 0;
        pixel_data[23][194] = 0;
        pixel_data[23][195] = 0;
        pixel_data[23][196] = 0;
        pixel_data[23][197] = 0;
        pixel_data[23][198] = 0;
        pixel_data[23][199] = 0; // y=23
        pixel_data[24][0] = 0;
        pixel_data[24][1] = 0;
        pixel_data[24][2] = 0;
        pixel_data[24][3] = 0;
        pixel_data[24][4] = 0;
        pixel_data[24][5] = 0;
        pixel_data[24][6] = 0;
        pixel_data[24][7] = 0;
        pixel_data[24][8] = 0;
        pixel_data[24][9] = 0;
        pixel_data[24][10] = 0;
        pixel_data[24][11] = 0;
        pixel_data[24][12] = 0;
        pixel_data[24][13] = 0;
        pixel_data[24][14] = 0;
        pixel_data[24][15] = 0;
        pixel_data[24][16] = 0;
        pixel_data[24][17] = 0;
        pixel_data[24][18] = 0;
        pixel_data[24][19] = 0;
        pixel_data[24][20] = 0;
        pixel_data[24][21] = 0;
        pixel_data[24][22] = 0;
        pixel_data[24][23] = 0;
        pixel_data[24][24] = 0;
        pixel_data[24][25] = 0;
        pixel_data[24][26] = 0;
        pixel_data[24][27] = 0;
        pixel_data[24][28] = 0;
        pixel_data[24][29] = 0;
        pixel_data[24][30] = 0;
        pixel_data[24][31] = 0;
        pixel_data[24][32] = 0;
        pixel_data[24][33] = 0;
        pixel_data[24][34] = 0;
        pixel_data[24][35] = 0;
        pixel_data[24][36] = 0;
        pixel_data[24][37] = 0;
        pixel_data[24][38] = 0;
        pixel_data[24][39] = 0;
        pixel_data[24][40] = 0;
        pixel_data[24][41] = 0;
        pixel_data[24][42] = 0;
        pixel_data[24][43] = 0;
        pixel_data[24][44] = 0;
        pixel_data[24][45] = 0;
        pixel_data[24][46] = 0;
        pixel_data[24][47] = 0;
        pixel_data[24][48] = 0;
        pixel_data[24][49] = 0;
        pixel_data[24][50] = 0;
        pixel_data[24][51] = 0;
        pixel_data[24][52] = 0;
        pixel_data[24][53] = 0;
        pixel_data[24][54] = 0;
        pixel_data[24][55] = 0;
        pixel_data[24][56] = 0;
        pixel_data[24][57] = 0;
        pixel_data[24][58] = 0;
        pixel_data[24][59] = 0;
        pixel_data[24][60] = 0;
        pixel_data[24][61] = 0;
        pixel_data[24][62] = 0;
        pixel_data[24][63] = 0;
        pixel_data[24][64] = 0;
        pixel_data[24][65] = 0;
        pixel_data[24][66] = 0;
        pixel_data[24][67] = 0;
        pixel_data[24][68] = 0;
        pixel_data[24][69] = 0;
        pixel_data[24][70] = 0;
        pixel_data[24][71] = 0;
        pixel_data[24][72] = 0;
        pixel_data[24][73] = 0;
        pixel_data[24][74] = 0;
        pixel_data[24][75] = 0;
        pixel_data[24][76] = 0;
        pixel_data[24][77] = 0;
        pixel_data[24][78] = 0;
        pixel_data[24][79] = 0;
        pixel_data[24][80] = 0;
        pixel_data[24][81] = 0;
        pixel_data[24][82] = 0;
        pixel_data[24][83] = 0;
        pixel_data[24][84] = 0;
        pixel_data[24][85] = 0;
        pixel_data[24][86] = 0;
        pixel_data[24][87] = 0;
        pixel_data[24][88] = 0;
        pixel_data[24][89] = 0;
        pixel_data[24][90] = 0;
        pixel_data[24][91] = 0;
        pixel_data[24][92] = 0;
        pixel_data[24][93] = 0;
        pixel_data[24][94] = 0;
        pixel_data[24][95] = 0;
        pixel_data[24][96] = 0;
        pixel_data[24][97] = 0;
        pixel_data[24][98] = 0;
        pixel_data[24][99] = 0;
        pixel_data[24][100] = 0;
        pixel_data[24][101] = 0;
        pixel_data[24][102] = 0;
        pixel_data[24][103] = 0;
        pixel_data[24][104] = 0;
        pixel_data[24][105] = 0;
        pixel_data[24][106] = 0;
        pixel_data[24][107] = 0;
        pixel_data[24][108] = 0;
        pixel_data[24][109] = 0;
        pixel_data[24][110] = 0;
        pixel_data[24][111] = 0;
        pixel_data[24][112] = 0;
        pixel_data[24][113] = 0;
        pixel_data[24][114] = 0;
        pixel_data[24][115] = 0;
        pixel_data[24][116] = 0;
        pixel_data[24][117] = 0;
        pixel_data[24][118] = 0;
        pixel_data[24][119] = 0;
        pixel_data[24][120] = 0;
        pixel_data[24][121] = 0;
        pixel_data[24][122] = 0;
        pixel_data[24][123] = 0;
        pixel_data[24][124] = 0;
        pixel_data[24][125] = 0;
        pixel_data[24][126] = 0;
        pixel_data[24][127] = 0;
        pixel_data[24][128] = 0;
        pixel_data[24][129] = 0;
        pixel_data[24][130] = 0;
        pixel_data[24][131] = 0;
        pixel_data[24][132] = 0;
        pixel_data[24][133] = 0;
        pixel_data[24][134] = 0;
        pixel_data[24][135] = 0;
        pixel_data[24][136] = 0;
        pixel_data[24][137] = 0;
        pixel_data[24][138] = 0;
        pixel_data[24][139] = 0;
        pixel_data[24][140] = 0;
        pixel_data[24][141] = 0;
        pixel_data[24][142] = 0;
        pixel_data[24][143] = 0;
        pixel_data[24][144] = 0;
        pixel_data[24][145] = 0;
        pixel_data[24][146] = 0;
        pixel_data[24][147] = 0;
        pixel_data[24][148] = 0;
        pixel_data[24][149] = 0;
        pixel_data[24][150] = 0;
        pixel_data[24][151] = 0;
        pixel_data[24][152] = 0;
        pixel_data[24][153] = 0;
        pixel_data[24][154] = 0;
        pixel_data[24][155] = 0;
        pixel_data[24][156] = 0;
        pixel_data[24][157] = 0;
        pixel_data[24][158] = 0;
        pixel_data[24][159] = 0;
        pixel_data[24][160] = 0;
        pixel_data[24][161] = 0;
        pixel_data[24][162] = 0;
        pixel_data[24][163] = 0;
        pixel_data[24][164] = 0;
        pixel_data[24][165] = 0;
        pixel_data[24][166] = 0;
        pixel_data[24][167] = 0;
        pixel_data[24][168] = 0;
        pixel_data[24][169] = 0;
        pixel_data[24][170] = 0;
        pixel_data[24][171] = 0;
        pixel_data[24][172] = 0;
        pixel_data[24][173] = 0;
        pixel_data[24][174] = 0;
        pixel_data[24][175] = 0;
        pixel_data[24][176] = 0;
        pixel_data[24][177] = 0;
        pixel_data[24][178] = 0;
        pixel_data[24][179] = 0;
        pixel_data[24][180] = 0;
        pixel_data[24][181] = 0;
        pixel_data[24][182] = 0;
        pixel_data[24][183] = 0;
        pixel_data[24][184] = 0;
        pixel_data[24][185] = 0;
        pixel_data[24][186] = 0;
        pixel_data[24][187] = 0;
        pixel_data[24][188] = 0;
        pixel_data[24][189] = 0;
        pixel_data[24][190] = 0;
        pixel_data[24][191] = 0;
        pixel_data[24][192] = 0;
        pixel_data[24][193] = 0;
        pixel_data[24][194] = 0;
        pixel_data[24][195] = 0;
        pixel_data[24][196] = 0;
        pixel_data[24][197] = 0;
        pixel_data[24][198] = 0;
        pixel_data[24][199] = 0; // y=24
        pixel_data[25][0] = 0;
        pixel_data[25][1] = 0;
        pixel_data[25][2] = 0;
        pixel_data[25][3] = 0;
        pixel_data[25][4] = 0;
        pixel_data[25][5] = 0;
        pixel_data[25][6] = 0;
        pixel_data[25][7] = 0;
        pixel_data[25][8] = 0;
        pixel_data[25][9] = 0;
        pixel_data[25][10] = 0;
        pixel_data[25][11] = 0;
        pixel_data[25][12] = 0;
        pixel_data[25][13] = 0;
        pixel_data[25][14] = 0;
        pixel_data[25][15] = 0;
        pixel_data[25][16] = 0;
        pixel_data[25][17] = 0;
        pixel_data[25][18] = 0;
        pixel_data[25][19] = 0;
        pixel_data[25][20] = 0;
        pixel_data[25][21] = 0;
        pixel_data[25][22] = 0;
        pixel_data[25][23] = 0;
        pixel_data[25][24] = 0;
        pixel_data[25][25] = 0;
        pixel_data[25][26] = 0;
        pixel_data[25][27] = 0;
        pixel_data[25][28] = 0;
        pixel_data[25][29] = 0;
        pixel_data[25][30] = 0;
        pixel_data[25][31] = 0;
        pixel_data[25][32] = 0;
        pixel_data[25][33] = 0;
        pixel_data[25][34] = 0;
        pixel_data[25][35] = 0;
        pixel_data[25][36] = 0;
        pixel_data[25][37] = 0;
        pixel_data[25][38] = 0;
        pixel_data[25][39] = 0;
        pixel_data[25][40] = 0;
        pixel_data[25][41] = 0;
        pixel_data[25][42] = 0;
        pixel_data[25][43] = 0;
        pixel_data[25][44] = 0;
        pixel_data[25][45] = 0;
        pixel_data[25][46] = 0;
        pixel_data[25][47] = 0;
        pixel_data[25][48] = 0;
        pixel_data[25][49] = 0;
        pixel_data[25][50] = 0;
        pixel_data[25][51] = 0;
        pixel_data[25][52] = 0;
        pixel_data[25][53] = 0;
        pixel_data[25][54] = 0;
        pixel_data[25][55] = 0;
        pixel_data[25][56] = 0;
        pixel_data[25][57] = 0;
        pixel_data[25][58] = 0;
        pixel_data[25][59] = 0;
        pixel_data[25][60] = 0;
        pixel_data[25][61] = 0;
        pixel_data[25][62] = 0;
        pixel_data[25][63] = 0;
        pixel_data[25][64] = 0;
        pixel_data[25][65] = 0;
        pixel_data[25][66] = 0;
        pixel_data[25][67] = 0;
        pixel_data[25][68] = 0;
        pixel_data[25][69] = 0;
        pixel_data[25][70] = 0;
        pixel_data[25][71] = 0;
        pixel_data[25][72] = 0;
        pixel_data[25][73] = 0;
        pixel_data[25][74] = 0;
        pixel_data[25][75] = 0;
        pixel_data[25][76] = 0;
        pixel_data[25][77] = 0;
        pixel_data[25][78] = 0;
        pixel_data[25][79] = 0;
        pixel_data[25][80] = 0;
        pixel_data[25][81] = 0;
        pixel_data[25][82] = 0;
        pixel_data[25][83] = 0;
        pixel_data[25][84] = 0;
        pixel_data[25][85] = 0;
        pixel_data[25][86] = 0;
        pixel_data[25][87] = 0;
        pixel_data[25][88] = 0;
        pixel_data[25][89] = 0;
        pixel_data[25][90] = 0;
        pixel_data[25][91] = 0;
        pixel_data[25][92] = 0;
        pixel_data[25][93] = 0;
        pixel_data[25][94] = 0;
        pixel_data[25][95] = 0;
        pixel_data[25][96] = 0;
        pixel_data[25][97] = 0;
        pixel_data[25][98] = 0;
        pixel_data[25][99] = 0;
        pixel_data[25][100] = 0;
        pixel_data[25][101] = 0;
        pixel_data[25][102] = 0;
        pixel_data[25][103] = 0;
        pixel_data[25][104] = 0;
        pixel_data[25][105] = 0;
        pixel_data[25][106] = 0;
        pixel_data[25][107] = 0;
        pixel_data[25][108] = 0;
        pixel_data[25][109] = 0;
        pixel_data[25][110] = 0;
        pixel_data[25][111] = 0;
        pixel_data[25][112] = 0;
        pixel_data[25][113] = 0;
        pixel_data[25][114] = 0;
        pixel_data[25][115] = 0;
        pixel_data[25][116] = 0;
        pixel_data[25][117] = 0;
        pixel_data[25][118] = 0;
        pixel_data[25][119] = 0;
        pixel_data[25][120] = 0;
        pixel_data[25][121] = 0;
        pixel_data[25][122] = 0;
        pixel_data[25][123] = 0;
        pixel_data[25][124] = 0;
        pixel_data[25][125] = 0;
        pixel_data[25][126] = 0;
        pixel_data[25][127] = 0;
        pixel_data[25][128] = 0;
        pixel_data[25][129] = 0;
        pixel_data[25][130] = 0;
        pixel_data[25][131] = 0;
        pixel_data[25][132] = 0;
        pixel_data[25][133] = 0;
        pixel_data[25][134] = 0;
        pixel_data[25][135] = 0;
        pixel_data[25][136] = 0;
        pixel_data[25][137] = 0;
        pixel_data[25][138] = 0;
        pixel_data[25][139] = 0;
        pixel_data[25][140] = 0;
        pixel_data[25][141] = 0;
        pixel_data[25][142] = 0;
        pixel_data[25][143] = 0;
        pixel_data[25][144] = 0;
        pixel_data[25][145] = 0;
        pixel_data[25][146] = 0;
        pixel_data[25][147] = 0;
        pixel_data[25][148] = 0;
        pixel_data[25][149] = 0;
        pixel_data[25][150] = 0;
        pixel_data[25][151] = 0;
        pixel_data[25][152] = 0;
        pixel_data[25][153] = 0;
        pixel_data[25][154] = 0;
        pixel_data[25][155] = 0;
        pixel_data[25][156] = 0;
        pixel_data[25][157] = 0;
        pixel_data[25][158] = 0;
        pixel_data[25][159] = 0;
        pixel_data[25][160] = 0;
        pixel_data[25][161] = 0;
        pixel_data[25][162] = 0;
        pixel_data[25][163] = 0;
        pixel_data[25][164] = 0;
        pixel_data[25][165] = 0;
        pixel_data[25][166] = 0;
        pixel_data[25][167] = 0;
        pixel_data[25][168] = 0;
        pixel_data[25][169] = 0;
        pixel_data[25][170] = 0;
        pixel_data[25][171] = 0;
        pixel_data[25][172] = 0;
        pixel_data[25][173] = 0;
        pixel_data[25][174] = 0;
        pixel_data[25][175] = 0;
        pixel_data[25][176] = 0;
        pixel_data[25][177] = 0;
        pixel_data[25][178] = 0;
        pixel_data[25][179] = 0;
        pixel_data[25][180] = 0;
        pixel_data[25][181] = 0;
        pixel_data[25][182] = 0;
        pixel_data[25][183] = 0;
        pixel_data[25][184] = 0;
        pixel_data[25][185] = 0;
        pixel_data[25][186] = 0;
        pixel_data[25][187] = 0;
        pixel_data[25][188] = 0;
        pixel_data[25][189] = 0;
        pixel_data[25][190] = 0;
        pixel_data[25][191] = 0;
        pixel_data[25][192] = 0;
        pixel_data[25][193] = 0;
        pixel_data[25][194] = 0;
        pixel_data[25][195] = 0;
        pixel_data[25][196] = 0;
        pixel_data[25][197] = 0;
        pixel_data[25][198] = 0;
        pixel_data[25][199] = 0; // y=25
        pixel_data[26][0] = 0;
        pixel_data[26][1] = 0;
        pixel_data[26][2] = 0;
        pixel_data[26][3] = 0;
        pixel_data[26][4] = 0;
        pixel_data[26][5] = 0;
        pixel_data[26][6] = 0;
        pixel_data[26][7] = 0;
        pixel_data[26][8] = 0;
        pixel_data[26][9] = 0;
        pixel_data[26][10] = 0;
        pixel_data[26][11] = 0;
        pixel_data[26][12] = 0;
        pixel_data[26][13] = 0;
        pixel_data[26][14] = 0;
        pixel_data[26][15] = 0;
        pixel_data[26][16] = 0;
        pixel_data[26][17] = 0;
        pixel_data[26][18] = 0;
        pixel_data[26][19] = 0;
        pixel_data[26][20] = 0;
        pixel_data[26][21] = 0;
        pixel_data[26][22] = 0;
        pixel_data[26][23] = 0;
        pixel_data[26][24] = 0;
        pixel_data[26][25] = 0;
        pixel_data[26][26] = 0;
        pixel_data[26][27] = 0;
        pixel_data[26][28] = 0;
        pixel_data[26][29] = 0;
        pixel_data[26][30] = 0;
        pixel_data[26][31] = 0;
        pixel_data[26][32] = 0;
        pixel_data[26][33] = 0;
        pixel_data[26][34] = 0;
        pixel_data[26][35] = 0;
        pixel_data[26][36] = 0;
        pixel_data[26][37] = 0;
        pixel_data[26][38] = 0;
        pixel_data[26][39] = 0;
        pixel_data[26][40] = 0;
        pixel_data[26][41] = 0;
        pixel_data[26][42] = 0;
        pixel_data[26][43] = 0;
        pixel_data[26][44] = 0;
        pixel_data[26][45] = 0;
        pixel_data[26][46] = 0;
        pixel_data[26][47] = 0;
        pixel_data[26][48] = 0;
        pixel_data[26][49] = 0;
        pixel_data[26][50] = 0;
        pixel_data[26][51] = 0;
        pixel_data[26][52] = 0;
        pixel_data[26][53] = 0;
        pixel_data[26][54] = 0;
        pixel_data[26][55] = 0;
        pixel_data[26][56] = 0;
        pixel_data[26][57] = 0;
        pixel_data[26][58] = 0;
        pixel_data[26][59] = 0;
        pixel_data[26][60] = 0;
        pixel_data[26][61] = 0;
        pixel_data[26][62] = 0;
        pixel_data[26][63] = 0;
        pixel_data[26][64] = 0;
        pixel_data[26][65] = 0;
        pixel_data[26][66] = 0;
        pixel_data[26][67] = 0;
        pixel_data[26][68] = 0;
        pixel_data[26][69] = 0;
        pixel_data[26][70] = 0;
        pixel_data[26][71] = 0;
        pixel_data[26][72] = 0;
        pixel_data[26][73] = 0;
        pixel_data[26][74] = 0;
        pixel_data[26][75] = 0;
        pixel_data[26][76] = 0;
        pixel_data[26][77] = 0;
        pixel_data[26][78] = 0;
        pixel_data[26][79] = 0;
        pixel_data[26][80] = 0;
        pixel_data[26][81] = 0;
        pixel_data[26][82] = 0;
        pixel_data[26][83] = 0;
        pixel_data[26][84] = 0;
        pixel_data[26][85] = 0;
        pixel_data[26][86] = 0;
        pixel_data[26][87] = 0;
        pixel_data[26][88] = 0;
        pixel_data[26][89] = 0;
        pixel_data[26][90] = 0;
        pixel_data[26][91] = 0;
        pixel_data[26][92] = 0;
        pixel_data[26][93] = 0;
        pixel_data[26][94] = 0;
        pixel_data[26][95] = 0;
        pixel_data[26][96] = 0;
        pixel_data[26][97] = 0;
        pixel_data[26][98] = 0;
        pixel_data[26][99] = 0;
        pixel_data[26][100] = 0;
        pixel_data[26][101] = 0;
        pixel_data[26][102] = 0;
        pixel_data[26][103] = 0;
        pixel_data[26][104] = 0;
        pixel_data[26][105] = 0;
        pixel_data[26][106] = 0;
        pixel_data[26][107] = 0;
        pixel_data[26][108] = 0;
        pixel_data[26][109] = 0;
        pixel_data[26][110] = 0;
        pixel_data[26][111] = 0;
        pixel_data[26][112] = 0;
        pixel_data[26][113] = 0;
        pixel_data[26][114] = 0;
        pixel_data[26][115] = 0;
        pixel_data[26][116] = 0;
        pixel_data[26][117] = 0;
        pixel_data[26][118] = 0;
        pixel_data[26][119] = 0;
        pixel_data[26][120] = 0;
        pixel_data[26][121] = 0;
        pixel_data[26][122] = 0;
        pixel_data[26][123] = 0;
        pixel_data[26][124] = 0;
        pixel_data[26][125] = 0;
        pixel_data[26][126] = 0;
        pixel_data[26][127] = 0;
        pixel_data[26][128] = 0;
        pixel_data[26][129] = 0;
        pixel_data[26][130] = 0;
        pixel_data[26][131] = 0;
        pixel_data[26][132] = 0;
        pixel_data[26][133] = 0;
        pixel_data[26][134] = 0;
        pixel_data[26][135] = 0;
        pixel_data[26][136] = 0;
        pixel_data[26][137] = 0;
        pixel_data[26][138] = 0;
        pixel_data[26][139] = 0;
        pixel_data[26][140] = 0;
        pixel_data[26][141] = 0;
        pixel_data[26][142] = 0;
        pixel_data[26][143] = 0;
        pixel_data[26][144] = 0;
        pixel_data[26][145] = 0;
        pixel_data[26][146] = 0;
        pixel_data[26][147] = 0;
        pixel_data[26][148] = 0;
        pixel_data[26][149] = 0;
        pixel_data[26][150] = 0;
        pixel_data[26][151] = 0;
        pixel_data[26][152] = 0;
        pixel_data[26][153] = 0;
        pixel_data[26][154] = 0;
        pixel_data[26][155] = 0;
        pixel_data[26][156] = 0;
        pixel_data[26][157] = 0;
        pixel_data[26][158] = 0;
        pixel_data[26][159] = 0;
        pixel_data[26][160] = 0;
        pixel_data[26][161] = 0;
        pixel_data[26][162] = 0;
        pixel_data[26][163] = 0;
        pixel_data[26][164] = 0;
        pixel_data[26][165] = 0;
        pixel_data[26][166] = 0;
        pixel_data[26][167] = 0;
        pixel_data[26][168] = 0;
        pixel_data[26][169] = 0;
        pixel_data[26][170] = 0;
        pixel_data[26][171] = 0;
        pixel_data[26][172] = 0;
        pixel_data[26][173] = 0;
        pixel_data[26][174] = 0;
        pixel_data[26][175] = 0;
        pixel_data[26][176] = 0;
        pixel_data[26][177] = 0;
        pixel_data[26][178] = 0;
        pixel_data[26][179] = 0;
        pixel_data[26][180] = 0;
        pixel_data[26][181] = 0;
        pixel_data[26][182] = 0;
        pixel_data[26][183] = 0;
        pixel_data[26][184] = 0;
        pixel_data[26][185] = 0;
        pixel_data[26][186] = 0;
        pixel_data[26][187] = 0;
        pixel_data[26][188] = 0;
        pixel_data[26][189] = 0;
        pixel_data[26][190] = 0;
        pixel_data[26][191] = 0;
        pixel_data[26][192] = 0;
        pixel_data[26][193] = 0;
        pixel_data[26][194] = 0;
        pixel_data[26][195] = 0;
        pixel_data[26][196] = 0;
        pixel_data[26][197] = 0;
        pixel_data[26][198] = 0;
        pixel_data[26][199] = 0; // y=26
        pixel_data[27][0] = 0;
        pixel_data[27][1] = 0;
        pixel_data[27][2] = 0;
        pixel_data[27][3] = 0;
        pixel_data[27][4] = 0;
        pixel_data[27][5] = 0;
        pixel_data[27][6] = 0;
        pixel_data[27][7] = 0;
        pixel_data[27][8] = 0;
        pixel_data[27][9] = 0;
        pixel_data[27][10] = 0;
        pixel_data[27][11] = 0;
        pixel_data[27][12] = 0;
        pixel_data[27][13] = 0;
        pixel_data[27][14] = 0;
        pixel_data[27][15] = 0;
        pixel_data[27][16] = 0;
        pixel_data[27][17] = 0;
        pixel_data[27][18] = 0;
        pixel_data[27][19] = 0;
        pixel_data[27][20] = 0;
        pixel_data[27][21] = 0;
        pixel_data[27][22] = 0;
        pixel_data[27][23] = 0;
        pixel_data[27][24] = 0;
        pixel_data[27][25] = 0;
        pixel_data[27][26] = 0;
        pixel_data[27][27] = 0;
        pixel_data[27][28] = 0;
        pixel_data[27][29] = 0;
        pixel_data[27][30] = 0;
        pixel_data[27][31] = 0;
        pixel_data[27][32] = 0;
        pixel_data[27][33] = 0;
        pixel_data[27][34] = 0;
        pixel_data[27][35] = 0;
        pixel_data[27][36] = 0;
        pixel_data[27][37] = 0;
        pixel_data[27][38] = 0;
        pixel_data[27][39] = 0;
        pixel_data[27][40] = 0;
        pixel_data[27][41] = 0;
        pixel_data[27][42] = 0;
        pixel_data[27][43] = 0;
        pixel_data[27][44] = 0;
        pixel_data[27][45] = 0;
        pixel_data[27][46] = 0;
        pixel_data[27][47] = 0;
        pixel_data[27][48] = 0;
        pixel_data[27][49] = 0;
        pixel_data[27][50] = 0;
        pixel_data[27][51] = 0;
        pixel_data[27][52] = 0;
        pixel_data[27][53] = 0;
        pixel_data[27][54] = 0;
        pixel_data[27][55] = 0;
        pixel_data[27][56] = 0;
        pixel_data[27][57] = 0;
        pixel_data[27][58] = 0;
        pixel_data[27][59] = 0;
        pixel_data[27][60] = 0;
        pixel_data[27][61] = 0;
        pixel_data[27][62] = 0;
        pixel_data[27][63] = 0;
        pixel_data[27][64] = 0;
        pixel_data[27][65] = 0;
        pixel_data[27][66] = 0;
        pixel_data[27][67] = 0;
        pixel_data[27][68] = 0;
        pixel_data[27][69] = 0;
        pixel_data[27][70] = 0;
        pixel_data[27][71] = 0;
        pixel_data[27][72] = 0;
        pixel_data[27][73] = 0;
        pixel_data[27][74] = 0;
        pixel_data[27][75] = 0;
        pixel_data[27][76] = 0;
        pixel_data[27][77] = 0;
        pixel_data[27][78] = 0;
        pixel_data[27][79] = 0;
        pixel_data[27][80] = 0;
        pixel_data[27][81] = 0;
        pixel_data[27][82] = 0;
        pixel_data[27][83] = 0;
        pixel_data[27][84] = 0;
        pixel_data[27][85] = 0;
        pixel_data[27][86] = 0;
        pixel_data[27][87] = 0;
        pixel_data[27][88] = 0;
        pixel_data[27][89] = 0;
        pixel_data[27][90] = 0;
        pixel_data[27][91] = 0;
        pixel_data[27][92] = 0;
        pixel_data[27][93] = 0;
        pixel_data[27][94] = 0;
        pixel_data[27][95] = 0;
        pixel_data[27][96] = 0;
        pixel_data[27][97] = 0;
        pixel_data[27][98] = 0;
        pixel_data[27][99] = 0;
        pixel_data[27][100] = 0;
        pixel_data[27][101] = 0;
        pixel_data[27][102] = 0;
        pixel_data[27][103] = 0;
        pixel_data[27][104] = 0;
        pixel_data[27][105] = 0;
        pixel_data[27][106] = 0;
        pixel_data[27][107] = 0;
        pixel_data[27][108] = 0;
        pixel_data[27][109] = 0;
        pixel_data[27][110] = 0;
        pixel_data[27][111] = 0;
        pixel_data[27][112] = 0;
        pixel_data[27][113] = 0;
        pixel_data[27][114] = 0;
        pixel_data[27][115] = 0;
        pixel_data[27][116] = 0;
        pixel_data[27][117] = 0;
        pixel_data[27][118] = 0;
        pixel_data[27][119] = 0;
        pixel_data[27][120] = 0;
        pixel_data[27][121] = 0;
        pixel_data[27][122] = 0;
        pixel_data[27][123] = 0;
        pixel_data[27][124] = 0;
        pixel_data[27][125] = 0;
        pixel_data[27][126] = 0;
        pixel_data[27][127] = 0;
        pixel_data[27][128] = 0;
        pixel_data[27][129] = 0;
        pixel_data[27][130] = 0;
        pixel_data[27][131] = 0;
        pixel_data[27][132] = 0;
        pixel_data[27][133] = 0;
        pixel_data[27][134] = 0;
        pixel_data[27][135] = 0;
        pixel_data[27][136] = 0;
        pixel_data[27][137] = 0;
        pixel_data[27][138] = 0;
        pixel_data[27][139] = 0;
        pixel_data[27][140] = 0;
        pixel_data[27][141] = 0;
        pixel_data[27][142] = 0;
        pixel_data[27][143] = 0;
        pixel_data[27][144] = 0;
        pixel_data[27][145] = 0;
        pixel_data[27][146] = 0;
        pixel_data[27][147] = 0;
        pixel_data[27][148] = 0;
        pixel_data[27][149] = 0;
        pixel_data[27][150] = 0;
        pixel_data[27][151] = 0;
        pixel_data[27][152] = 0;
        pixel_data[27][153] = 0;
        pixel_data[27][154] = 0;
        pixel_data[27][155] = 0;
        pixel_data[27][156] = 0;
        pixel_data[27][157] = 0;
        pixel_data[27][158] = 0;
        pixel_data[27][159] = 0;
        pixel_data[27][160] = 0;
        pixel_data[27][161] = 0;
        pixel_data[27][162] = 0;
        pixel_data[27][163] = 0;
        pixel_data[27][164] = 0;
        pixel_data[27][165] = 0;
        pixel_data[27][166] = 0;
        pixel_data[27][167] = 0;
        pixel_data[27][168] = 0;
        pixel_data[27][169] = 0;
        pixel_data[27][170] = 0;
        pixel_data[27][171] = 0;
        pixel_data[27][172] = 0;
        pixel_data[27][173] = 0;
        pixel_data[27][174] = 0;
        pixel_data[27][175] = 0;
        pixel_data[27][176] = 0;
        pixel_data[27][177] = 0;
        pixel_data[27][178] = 0;
        pixel_data[27][179] = 0;
        pixel_data[27][180] = 0;
        pixel_data[27][181] = 0;
        pixel_data[27][182] = 0;
        pixel_data[27][183] = 0;
        pixel_data[27][184] = 0;
        pixel_data[27][185] = 0;
        pixel_data[27][186] = 0;
        pixel_data[27][187] = 0;
        pixel_data[27][188] = 0;
        pixel_data[27][189] = 0;
        pixel_data[27][190] = 0;
        pixel_data[27][191] = 0;
        pixel_data[27][192] = 0;
        pixel_data[27][193] = 0;
        pixel_data[27][194] = 0;
        pixel_data[27][195] = 0;
        pixel_data[27][196] = 0;
        pixel_data[27][197] = 0;
        pixel_data[27][198] = 0;
        pixel_data[27][199] = 0; // y=27
        pixel_data[28][0] = 0;
        pixel_data[28][1] = 0;
        pixel_data[28][2] = 0;
        pixel_data[28][3] = 0;
        pixel_data[28][4] = 0;
        pixel_data[28][5] = 0;
        pixel_data[28][6] = 0;
        pixel_data[28][7] = 0;
        pixel_data[28][8] = 0;
        pixel_data[28][9] = 0;
        pixel_data[28][10] = 0;
        pixel_data[28][11] = 0;
        pixel_data[28][12] = 0;
        pixel_data[28][13] = 0;
        pixel_data[28][14] = 0;
        pixel_data[28][15] = 0;
        pixel_data[28][16] = 0;
        pixel_data[28][17] = 0;
        pixel_data[28][18] = 0;
        pixel_data[28][19] = 0;
        pixel_data[28][20] = 0;
        pixel_data[28][21] = 0;
        pixel_data[28][22] = 0;
        pixel_data[28][23] = 0;
        pixel_data[28][24] = 0;
        pixel_data[28][25] = 0;
        pixel_data[28][26] = 0;
        pixel_data[28][27] = 0;
        pixel_data[28][28] = 0;
        pixel_data[28][29] = 0;
        pixel_data[28][30] = 0;
        pixel_data[28][31] = 0;
        pixel_data[28][32] = 0;
        pixel_data[28][33] = 0;
        pixel_data[28][34] = 0;
        pixel_data[28][35] = 0;
        pixel_data[28][36] = 0;
        pixel_data[28][37] = 0;
        pixel_data[28][38] = 0;
        pixel_data[28][39] = 0;
        pixel_data[28][40] = 0;
        pixel_data[28][41] = 0;
        pixel_data[28][42] = 0;
        pixel_data[28][43] = 0;
        pixel_data[28][44] = 0;
        pixel_data[28][45] = 0;
        pixel_data[28][46] = 0;
        pixel_data[28][47] = 0;
        pixel_data[28][48] = 0;
        pixel_data[28][49] = 0;
        pixel_data[28][50] = 0;
        pixel_data[28][51] = 0;
        pixel_data[28][52] = 0;
        pixel_data[28][53] = 0;
        pixel_data[28][54] = 0;
        pixel_data[28][55] = 0;
        pixel_data[28][56] = 0;
        pixel_data[28][57] = 0;
        pixel_data[28][58] = 0;
        pixel_data[28][59] = 0;
        pixel_data[28][60] = 0;
        pixel_data[28][61] = 0;
        pixel_data[28][62] = 0;
        pixel_data[28][63] = 0;
        pixel_data[28][64] = 0;
        pixel_data[28][65] = 0;
        pixel_data[28][66] = 0;
        pixel_data[28][67] = 0;
        pixel_data[28][68] = 0;
        pixel_data[28][69] = 0;
        pixel_data[28][70] = 0;
        pixel_data[28][71] = 0;
        pixel_data[28][72] = 0;
        pixel_data[28][73] = 0;
        pixel_data[28][74] = 0;
        pixel_data[28][75] = 0;
        pixel_data[28][76] = 0;
        pixel_data[28][77] = 0;
        pixel_data[28][78] = 0;
        pixel_data[28][79] = 0;
        pixel_data[28][80] = 0;
        pixel_data[28][81] = 0;
        pixel_data[28][82] = 0;
        pixel_data[28][83] = 0;
        pixel_data[28][84] = 0;
        pixel_data[28][85] = 0;
        pixel_data[28][86] = 0;
        pixel_data[28][87] = 0;
        pixel_data[28][88] = 0;
        pixel_data[28][89] = 0;
        pixel_data[28][90] = 0;
        pixel_data[28][91] = 0;
        pixel_data[28][92] = 0;
        pixel_data[28][93] = 0;
        pixel_data[28][94] = 0;
        pixel_data[28][95] = 0;
        pixel_data[28][96] = 0;
        pixel_data[28][97] = 0;
        pixel_data[28][98] = 0;
        pixel_data[28][99] = 0;
        pixel_data[28][100] = 0;
        pixel_data[28][101] = 0;
        pixel_data[28][102] = 0;
        pixel_data[28][103] = 0;
        pixel_data[28][104] = 0;
        pixel_data[28][105] = 0;
        pixel_data[28][106] = 0;
        pixel_data[28][107] = 0;
        pixel_data[28][108] = 0;
        pixel_data[28][109] = 0;
        pixel_data[28][110] = 0;
        pixel_data[28][111] = 0;
        pixel_data[28][112] = 0;
        pixel_data[28][113] = 0;
        pixel_data[28][114] = 0;
        pixel_data[28][115] = 0;
        pixel_data[28][116] = 0;
        pixel_data[28][117] = 0;
        pixel_data[28][118] = 0;
        pixel_data[28][119] = 0;
        pixel_data[28][120] = 0;
        pixel_data[28][121] = 0;
        pixel_data[28][122] = 0;
        pixel_data[28][123] = 0;
        pixel_data[28][124] = 0;
        pixel_data[28][125] = 0;
        pixel_data[28][126] = 0;
        pixel_data[28][127] = 0;
        pixel_data[28][128] = 0;
        pixel_data[28][129] = 0;
        pixel_data[28][130] = 0;
        pixel_data[28][131] = 0;
        pixel_data[28][132] = 0;
        pixel_data[28][133] = 0;
        pixel_data[28][134] = 0;
        pixel_data[28][135] = 0;
        pixel_data[28][136] = 0;
        pixel_data[28][137] = 0;
        pixel_data[28][138] = 0;
        pixel_data[28][139] = 0;
        pixel_data[28][140] = 0;
        pixel_data[28][141] = 0;
        pixel_data[28][142] = 0;
        pixel_data[28][143] = 0;
        pixel_data[28][144] = 0;
        pixel_data[28][145] = 0;
        pixel_data[28][146] = 0;
        pixel_data[28][147] = 0;
        pixel_data[28][148] = 0;
        pixel_data[28][149] = 0;
        pixel_data[28][150] = 0;
        pixel_data[28][151] = 0;
        pixel_data[28][152] = 0;
        pixel_data[28][153] = 0;
        pixel_data[28][154] = 0;
        pixel_data[28][155] = 0;
        pixel_data[28][156] = 0;
        pixel_data[28][157] = 0;
        pixel_data[28][158] = 0;
        pixel_data[28][159] = 0;
        pixel_data[28][160] = 0;
        pixel_data[28][161] = 0;
        pixel_data[28][162] = 0;
        pixel_data[28][163] = 0;
        pixel_data[28][164] = 0;
        pixel_data[28][165] = 0;
        pixel_data[28][166] = 0;
        pixel_data[28][167] = 0;
        pixel_data[28][168] = 0;
        pixel_data[28][169] = 0;
        pixel_data[28][170] = 0;
        pixel_data[28][171] = 0;
        pixel_data[28][172] = 0;
        pixel_data[28][173] = 0;
        pixel_data[28][174] = 0;
        pixel_data[28][175] = 0;
        pixel_data[28][176] = 0;
        pixel_data[28][177] = 0;
        pixel_data[28][178] = 0;
        pixel_data[28][179] = 0;
        pixel_data[28][180] = 0;
        pixel_data[28][181] = 0;
        pixel_data[28][182] = 0;
        pixel_data[28][183] = 0;
        pixel_data[28][184] = 0;
        pixel_data[28][185] = 0;
        pixel_data[28][186] = 0;
        pixel_data[28][187] = 0;
        pixel_data[28][188] = 0;
        pixel_data[28][189] = 0;
        pixel_data[28][190] = 0;
        pixel_data[28][191] = 0;
        pixel_data[28][192] = 0;
        pixel_data[28][193] = 0;
        pixel_data[28][194] = 0;
        pixel_data[28][195] = 0;
        pixel_data[28][196] = 0;
        pixel_data[28][197] = 0;
        pixel_data[28][198] = 0;
        pixel_data[28][199] = 0; // y=28
        pixel_data[29][0] = 0;
        pixel_data[29][1] = 0;
        pixel_data[29][2] = 0;
        pixel_data[29][3] = 0;
        pixel_data[29][4] = 0;
        pixel_data[29][5] = 0;
        pixel_data[29][6] = 0;
        pixel_data[29][7] = 0;
        pixel_data[29][8] = 0;
        pixel_data[29][9] = 0;
        pixel_data[29][10] = 0;
        pixel_data[29][11] = 0;
        pixel_data[29][12] = 0;
        pixel_data[29][13] = 0;
        pixel_data[29][14] = 0;
        pixel_data[29][15] = 0;
        pixel_data[29][16] = 0;
        pixel_data[29][17] = 0;
        pixel_data[29][18] = 0;
        pixel_data[29][19] = 0;
        pixel_data[29][20] = 0;
        pixel_data[29][21] = 0;
        pixel_data[29][22] = 0;
        pixel_data[29][23] = 0;
        pixel_data[29][24] = 0;
        pixel_data[29][25] = 0;
        pixel_data[29][26] = 0;
        pixel_data[29][27] = 0;
        pixel_data[29][28] = 0;
        pixel_data[29][29] = 0;
        pixel_data[29][30] = 0;
        pixel_data[29][31] = 0;
        pixel_data[29][32] = 0;
        pixel_data[29][33] = 0;
        pixel_data[29][34] = 0;
        pixel_data[29][35] = 0;
        pixel_data[29][36] = 0;
        pixel_data[29][37] = 0;
        pixel_data[29][38] = 0;
        pixel_data[29][39] = 0;
        pixel_data[29][40] = 0;
        pixel_data[29][41] = 0;
        pixel_data[29][42] = 0;
        pixel_data[29][43] = 0;
        pixel_data[29][44] = 0;
        pixel_data[29][45] = 0;
        pixel_data[29][46] = 0;
        pixel_data[29][47] = 0;
        pixel_data[29][48] = 0;
        pixel_data[29][49] = 0;
        pixel_data[29][50] = 0;
        pixel_data[29][51] = 0;
        pixel_data[29][52] = 0;
        pixel_data[29][53] = 0;
        pixel_data[29][54] = 0;
        pixel_data[29][55] = 0;
        pixel_data[29][56] = 0;
        pixel_data[29][57] = 0;
        pixel_data[29][58] = 0;
        pixel_data[29][59] = 0;
        pixel_data[29][60] = 0;
        pixel_data[29][61] = 0;
        pixel_data[29][62] = 0;
        pixel_data[29][63] = 0;
        pixel_data[29][64] = 0;
        pixel_data[29][65] = 0;
        pixel_data[29][66] = 0;
        pixel_data[29][67] = 0;
        pixel_data[29][68] = 0;
        pixel_data[29][69] = 0;
        pixel_data[29][70] = 0;
        pixel_data[29][71] = 0;
        pixel_data[29][72] = 0;
        pixel_data[29][73] = 0;
        pixel_data[29][74] = 0;
        pixel_data[29][75] = 0;
        pixel_data[29][76] = 0;
        pixel_data[29][77] = 0;
        pixel_data[29][78] = 0;
        pixel_data[29][79] = 0;
        pixel_data[29][80] = 0;
        pixel_data[29][81] = 0;
        pixel_data[29][82] = 0;
        pixel_data[29][83] = 0;
        pixel_data[29][84] = 0;
        pixel_data[29][85] = 0;
        pixel_data[29][86] = 0;
        pixel_data[29][87] = 0;
        pixel_data[29][88] = 0;
        pixel_data[29][89] = 0;
        pixel_data[29][90] = 0;
        pixel_data[29][91] = 0;
        pixel_data[29][92] = 0;
        pixel_data[29][93] = 0;
        pixel_data[29][94] = 0;
        pixel_data[29][95] = 0;
        pixel_data[29][96] = 0;
        pixel_data[29][97] = 0;
        pixel_data[29][98] = 0;
        pixel_data[29][99] = 0;
        pixel_data[29][100] = 0;
        pixel_data[29][101] = 0;
        pixel_data[29][102] = 0;
        pixel_data[29][103] = 0;
        pixel_data[29][104] = 0;
        pixel_data[29][105] = 0;
        pixel_data[29][106] = 0;
        pixel_data[29][107] = 0;
        pixel_data[29][108] = 0;
        pixel_data[29][109] = 0;
        pixel_data[29][110] = 0;
        pixel_data[29][111] = 0;
        pixel_data[29][112] = 0;
        pixel_data[29][113] = 0;
        pixel_data[29][114] = 0;
        pixel_data[29][115] = 0;
        pixel_data[29][116] = 0;
        pixel_data[29][117] = 0;
        pixel_data[29][118] = 0;
        pixel_data[29][119] = 0;
        pixel_data[29][120] = 0;
        pixel_data[29][121] = 0;
        pixel_data[29][122] = 0;
        pixel_data[29][123] = 0;
        pixel_data[29][124] = 0;
        pixel_data[29][125] = 0;
        pixel_data[29][126] = 0;
        pixel_data[29][127] = 0;
        pixel_data[29][128] = 0;
        pixel_data[29][129] = 0;
        pixel_data[29][130] = 0;
        pixel_data[29][131] = 0;
        pixel_data[29][132] = 0;
        pixel_data[29][133] = 0;
        pixel_data[29][134] = 0;
        pixel_data[29][135] = 0;
        pixel_data[29][136] = 0;
        pixel_data[29][137] = 0;
        pixel_data[29][138] = 0;
        pixel_data[29][139] = 0;
        pixel_data[29][140] = 0;
        pixel_data[29][141] = 0;
        pixel_data[29][142] = 0;
        pixel_data[29][143] = 0;
        pixel_data[29][144] = 0;
        pixel_data[29][145] = 0;
        pixel_data[29][146] = 0;
        pixel_data[29][147] = 0;
        pixel_data[29][148] = 0;
        pixel_data[29][149] = 0;
        pixel_data[29][150] = 0;
        pixel_data[29][151] = 0;
        pixel_data[29][152] = 0;
        pixel_data[29][153] = 0;
        pixel_data[29][154] = 0;
        pixel_data[29][155] = 0;
        pixel_data[29][156] = 0;
        pixel_data[29][157] = 0;
        pixel_data[29][158] = 0;
        pixel_data[29][159] = 0;
        pixel_data[29][160] = 0;
        pixel_data[29][161] = 0;
        pixel_data[29][162] = 0;
        pixel_data[29][163] = 0;
        pixel_data[29][164] = 0;
        pixel_data[29][165] = 0;
        pixel_data[29][166] = 0;
        pixel_data[29][167] = 0;
        pixel_data[29][168] = 0;
        pixel_data[29][169] = 0;
        pixel_data[29][170] = 0;
        pixel_data[29][171] = 0;
        pixel_data[29][172] = 0;
        pixel_data[29][173] = 0;
        pixel_data[29][174] = 0;
        pixel_data[29][175] = 0;
        pixel_data[29][176] = 0;
        pixel_data[29][177] = 0;
        pixel_data[29][178] = 0;
        pixel_data[29][179] = 0;
        pixel_data[29][180] = 0;
        pixel_data[29][181] = 0;
        pixel_data[29][182] = 0;
        pixel_data[29][183] = 0;
        pixel_data[29][184] = 0;
        pixel_data[29][185] = 0;
        pixel_data[29][186] = 0;
        pixel_data[29][187] = 0;
        pixel_data[29][188] = 0;
        pixel_data[29][189] = 0;
        pixel_data[29][190] = 0;
        pixel_data[29][191] = 0;
        pixel_data[29][192] = 0;
        pixel_data[29][193] = 0;
        pixel_data[29][194] = 0;
        pixel_data[29][195] = 0;
        pixel_data[29][196] = 0;
        pixel_data[29][197] = 0;
        pixel_data[29][198] = 0;
        pixel_data[29][199] = 0; // y=29
        pixel_data[30][0] = 0;
        pixel_data[30][1] = 0;
        pixel_data[30][2] = 0;
        pixel_data[30][3] = 0;
        pixel_data[30][4] = 0;
        pixel_data[30][5] = 0;
        pixel_data[30][6] = 0;
        pixel_data[30][7] = 0;
        pixel_data[30][8] = 0;
        pixel_data[30][9] = 0;
        pixel_data[30][10] = 0;
        pixel_data[30][11] = 0;
        pixel_data[30][12] = 0;
        pixel_data[30][13] = 0;
        pixel_data[30][14] = 0;
        pixel_data[30][15] = 0;
        pixel_data[30][16] = 0;
        pixel_data[30][17] = 0;
        pixel_data[30][18] = 0;
        pixel_data[30][19] = 0;
        pixel_data[30][20] = 0;
        pixel_data[30][21] = 0;
        pixel_data[30][22] = 0;
        pixel_data[30][23] = 0;
        pixel_data[30][24] = 0;
        pixel_data[30][25] = 0;
        pixel_data[30][26] = 0;
        pixel_data[30][27] = 0;
        pixel_data[30][28] = 0;
        pixel_data[30][29] = 0;
        pixel_data[30][30] = 0;
        pixel_data[30][31] = 0;
        pixel_data[30][32] = 0;
        pixel_data[30][33] = 0;
        pixel_data[30][34] = 0;
        pixel_data[30][35] = 0;
        pixel_data[30][36] = 0;
        pixel_data[30][37] = 0;
        pixel_data[30][38] = 0;
        pixel_data[30][39] = 0;
        pixel_data[30][40] = 0;
        pixel_data[30][41] = 0;
        pixel_data[30][42] = 0;
        pixel_data[30][43] = 0;
        pixel_data[30][44] = 0;
        pixel_data[30][45] = 0;
        pixel_data[30][46] = 0;
        pixel_data[30][47] = 0;
        pixel_data[30][48] = 0;
        pixel_data[30][49] = 0;
        pixel_data[30][50] = 0;
        pixel_data[30][51] = 0;
        pixel_data[30][52] = 0;
        pixel_data[30][53] = 0;
        pixel_data[30][54] = 0;
        pixel_data[30][55] = 0;
        pixel_data[30][56] = 0;
        pixel_data[30][57] = 0;
        pixel_data[30][58] = 0;
        pixel_data[30][59] = 0;
        pixel_data[30][60] = 0;
        pixel_data[30][61] = 0;
        pixel_data[30][62] = 0;
        pixel_data[30][63] = 0;
        pixel_data[30][64] = 0;
        pixel_data[30][65] = 0;
        pixel_data[30][66] = 0;
        pixel_data[30][67] = 0;
        pixel_data[30][68] = 0;
        pixel_data[30][69] = 0;
        pixel_data[30][70] = 0;
        pixel_data[30][71] = 0;
        pixel_data[30][72] = 0;
        pixel_data[30][73] = 0;
        pixel_data[30][74] = 0;
        pixel_data[30][75] = 0;
        pixel_data[30][76] = 0;
        pixel_data[30][77] = 0;
        pixel_data[30][78] = 0;
        pixel_data[30][79] = 0;
        pixel_data[30][80] = 0;
        pixel_data[30][81] = 0;
        pixel_data[30][82] = 0;
        pixel_data[30][83] = 0;
        pixel_data[30][84] = 0;
        pixel_data[30][85] = 0;
        pixel_data[30][86] = 0;
        pixel_data[30][87] = 0;
        pixel_data[30][88] = 0;
        pixel_data[30][89] = 0;
        pixel_data[30][90] = 0;
        pixel_data[30][91] = 0;
        pixel_data[30][92] = 0;
        pixel_data[30][93] = 0;
        pixel_data[30][94] = 0;
        pixel_data[30][95] = 0;
        pixel_data[30][96] = 0;
        pixel_data[30][97] = 0;
        pixel_data[30][98] = 0;
        pixel_data[30][99] = 0;
        pixel_data[30][100] = 0;
        pixel_data[30][101] = 0;
        pixel_data[30][102] = 0;
        pixel_data[30][103] = 0;
        pixel_data[30][104] = 0;
        pixel_data[30][105] = 0;
        pixel_data[30][106] = 0;
        pixel_data[30][107] = 0;
        pixel_data[30][108] = 0;
        pixel_data[30][109] = 0;
        pixel_data[30][110] = 0;
        pixel_data[30][111] = 0;
        pixel_data[30][112] = 0;
        pixel_data[30][113] = 0;
        pixel_data[30][114] = 0;
        pixel_data[30][115] = 0;
        pixel_data[30][116] = 0;
        pixel_data[30][117] = 0;
        pixel_data[30][118] = 0;
        pixel_data[30][119] = 0;
        pixel_data[30][120] = 0;
        pixel_data[30][121] = 0;
        pixel_data[30][122] = 0;
        pixel_data[30][123] = 0;
        pixel_data[30][124] = 0;
        pixel_data[30][125] = 0;
        pixel_data[30][126] = 0;
        pixel_data[30][127] = 0;
        pixel_data[30][128] = 0;
        pixel_data[30][129] = 0;
        pixel_data[30][130] = 0;
        pixel_data[30][131] = 0;
        pixel_data[30][132] = 0;
        pixel_data[30][133] = 0;
        pixel_data[30][134] = 0;
        pixel_data[30][135] = 0;
        pixel_data[30][136] = 0;
        pixel_data[30][137] = 0;
        pixel_data[30][138] = 0;
        pixel_data[30][139] = 0;
        pixel_data[30][140] = 0;
        pixel_data[30][141] = 0;
        pixel_data[30][142] = 0;
        pixel_data[30][143] = 0;
        pixel_data[30][144] = 0;
        pixel_data[30][145] = 0;
        pixel_data[30][146] = 0;
        pixel_data[30][147] = 0;
        pixel_data[30][148] = 0;
        pixel_data[30][149] = 0;
        pixel_data[30][150] = 0;
        pixel_data[30][151] = 0;
        pixel_data[30][152] = 0;
        pixel_data[30][153] = 0;
        pixel_data[30][154] = 0;
        pixel_data[30][155] = 0;
        pixel_data[30][156] = 0;
        pixel_data[30][157] = 0;
        pixel_data[30][158] = 0;
        pixel_data[30][159] = 0;
        pixel_data[30][160] = 0;
        pixel_data[30][161] = 0;
        pixel_data[30][162] = 0;
        pixel_data[30][163] = 0;
        pixel_data[30][164] = 0;
        pixel_data[30][165] = 0;
        pixel_data[30][166] = 0;
        pixel_data[30][167] = 0;
        pixel_data[30][168] = 0;
        pixel_data[30][169] = 0;
        pixel_data[30][170] = 0;
        pixel_data[30][171] = 0;
        pixel_data[30][172] = 0;
        pixel_data[30][173] = 0;
        pixel_data[30][174] = 0;
        pixel_data[30][175] = 0;
        pixel_data[30][176] = 0;
        pixel_data[30][177] = 0;
        pixel_data[30][178] = 0;
        pixel_data[30][179] = 0;
        pixel_data[30][180] = 0;
        pixel_data[30][181] = 0;
        pixel_data[30][182] = 0;
        pixel_data[30][183] = 0;
        pixel_data[30][184] = 0;
        pixel_data[30][185] = 0;
        pixel_data[30][186] = 0;
        pixel_data[30][187] = 0;
        pixel_data[30][188] = 0;
        pixel_data[30][189] = 0;
        pixel_data[30][190] = 0;
        pixel_data[30][191] = 0;
        pixel_data[30][192] = 0;
        pixel_data[30][193] = 0;
        pixel_data[30][194] = 0;
        pixel_data[30][195] = 0;
        pixel_data[30][196] = 0;
        pixel_data[30][197] = 0;
        pixel_data[30][198] = 0;
        pixel_data[30][199] = 0; // y=30
        pixel_data[31][0] = 0;
        pixel_data[31][1] = 0;
        pixel_data[31][2] = 0;
        pixel_data[31][3] = 0;
        pixel_data[31][4] = 0;
        pixel_data[31][5] = 0;
        pixel_data[31][6] = 0;
        pixel_data[31][7] = 0;
        pixel_data[31][8] = 0;
        pixel_data[31][9] = 0;
        pixel_data[31][10] = 0;
        pixel_data[31][11] = 0;
        pixel_data[31][12] = 0;
        pixel_data[31][13] = 0;
        pixel_data[31][14] = 0;
        pixel_data[31][15] = 0;
        pixel_data[31][16] = 0;
        pixel_data[31][17] = 0;
        pixel_data[31][18] = 0;
        pixel_data[31][19] = 0;
        pixel_data[31][20] = 0;
        pixel_data[31][21] = 0;
        pixel_data[31][22] = 0;
        pixel_data[31][23] = 0;
        pixel_data[31][24] = 0;
        pixel_data[31][25] = 0;
        pixel_data[31][26] = 0;
        pixel_data[31][27] = 0;
        pixel_data[31][28] = 0;
        pixel_data[31][29] = 0;
        pixel_data[31][30] = 0;
        pixel_data[31][31] = 0;
        pixel_data[31][32] = 0;
        pixel_data[31][33] = 0;
        pixel_data[31][34] = 0;
        pixel_data[31][35] = 0;
        pixel_data[31][36] = 0;
        pixel_data[31][37] = 0;
        pixel_data[31][38] = 0;
        pixel_data[31][39] = 0;
        pixel_data[31][40] = 0;
        pixel_data[31][41] = 0;
        pixel_data[31][42] = 0;
        pixel_data[31][43] = 0;
        pixel_data[31][44] = 0;
        pixel_data[31][45] = 0;
        pixel_data[31][46] = 0;
        pixel_data[31][47] = 0;
        pixel_data[31][48] = 0;
        pixel_data[31][49] = 0;
        pixel_data[31][50] = 0;
        pixel_data[31][51] = 0;
        pixel_data[31][52] = 0;
        pixel_data[31][53] = 0;
        pixel_data[31][54] = 0;
        pixel_data[31][55] = 0;
        pixel_data[31][56] = 0;
        pixel_data[31][57] = 0;
        pixel_data[31][58] = 0;
        pixel_data[31][59] = 0;
        pixel_data[31][60] = 0;
        pixel_data[31][61] = 0;
        pixel_data[31][62] = 0;
        pixel_data[31][63] = 0;
        pixel_data[31][64] = 0;
        pixel_data[31][65] = 0;
        pixel_data[31][66] = 0;
        pixel_data[31][67] = 0;
        pixel_data[31][68] = 0;
        pixel_data[31][69] = 0;
        pixel_data[31][70] = 0;
        pixel_data[31][71] = 0;
        pixel_data[31][72] = 0;
        pixel_data[31][73] = 0;
        pixel_data[31][74] = 0;
        pixel_data[31][75] = 0;
        pixel_data[31][76] = 0;
        pixel_data[31][77] = 0;
        pixel_data[31][78] = 0;
        pixel_data[31][79] = 0;
        pixel_data[31][80] = 0;
        pixel_data[31][81] = 0;
        pixel_data[31][82] = 0;
        pixel_data[31][83] = 0;
        pixel_data[31][84] = 0;
        pixel_data[31][85] = 0;
        pixel_data[31][86] = 0;
        pixel_data[31][87] = 0;
        pixel_data[31][88] = 0;
        pixel_data[31][89] = 0;
        pixel_data[31][90] = 0;
        pixel_data[31][91] = 0;
        pixel_data[31][92] = 0;
        pixel_data[31][93] = 0;
        pixel_data[31][94] = 0;
        pixel_data[31][95] = 0;
        pixel_data[31][96] = 0;
        pixel_data[31][97] = 0;
        pixel_data[31][98] = 0;
        pixel_data[31][99] = 0;
        pixel_data[31][100] = 0;
        pixel_data[31][101] = 0;
        pixel_data[31][102] = 0;
        pixel_data[31][103] = 0;
        pixel_data[31][104] = 0;
        pixel_data[31][105] = 0;
        pixel_data[31][106] = 0;
        pixel_data[31][107] = 0;
        pixel_data[31][108] = 0;
        pixel_data[31][109] = 0;
        pixel_data[31][110] = 0;
        pixel_data[31][111] = 0;
        pixel_data[31][112] = 0;
        pixel_data[31][113] = 0;
        pixel_data[31][114] = 0;
        pixel_data[31][115] = 0;
        pixel_data[31][116] = 0;
        pixel_data[31][117] = 0;
        pixel_data[31][118] = 0;
        pixel_data[31][119] = 0;
        pixel_data[31][120] = 0;
        pixel_data[31][121] = 0;
        pixel_data[31][122] = 0;
        pixel_data[31][123] = 0;
        pixel_data[31][124] = 0;
        pixel_data[31][125] = 0;
        pixel_data[31][126] = 0;
        pixel_data[31][127] = 0;
        pixel_data[31][128] = 0;
        pixel_data[31][129] = 0;
        pixel_data[31][130] = 0;
        pixel_data[31][131] = 0;
        pixel_data[31][132] = 0;
        pixel_data[31][133] = 0;
        pixel_data[31][134] = 0;
        pixel_data[31][135] = 0;
        pixel_data[31][136] = 0;
        pixel_data[31][137] = 0;
        pixel_data[31][138] = 0;
        pixel_data[31][139] = 0;
        pixel_data[31][140] = 0;
        pixel_data[31][141] = 0;
        pixel_data[31][142] = 0;
        pixel_data[31][143] = 0;
        pixel_data[31][144] = 0;
        pixel_data[31][145] = 0;
        pixel_data[31][146] = 0;
        pixel_data[31][147] = 0;
        pixel_data[31][148] = 0;
        pixel_data[31][149] = 0;
        pixel_data[31][150] = 0;
        pixel_data[31][151] = 0;
        pixel_data[31][152] = 0;
        pixel_data[31][153] = 0;
        pixel_data[31][154] = 0;
        pixel_data[31][155] = 0;
        pixel_data[31][156] = 0;
        pixel_data[31][157] = 0;
        pixel_data[31][158] = 0;
        pixel_data[31][159] = 0;
        pixel_data[31][160] = 0;
        pixel_data[31][161] = 0;
        pixel_data[31][162] = 0;
        pixel_data[31][163] = 0;
        pixel_data[31][164] = 0;
        pixel_data[31][165] = 0;
        pixel_data[31][166] = 0;
        pixel_data[31][167] = 0;
        pixel_data[31][168] = 0;
        pixel_data[31][169] = 0;
        pixel_data[31][170] = 0;
        pixel_data[31][171] = 0;
        pixel_data[31][172] = 0;
        pixel_data[31][173] = 0;
        pixel_data[31][174] = 0;
        pixel_data[31][175] = 0;
        pixel_data[31][176] = 0;
        pixel_data[31][177] = 0;
        pixel_data[31][178] = 0;
        pixel_data[31][179] = 0;
        pixel_data[31][180] = 0;
        pixel_data[31][181] = 0;
        pixel_data[31][182] = 0;
        pixel_data[31][183] = 0;
        pixel_data[31][184] = 0;
        pixel_data[31][185] = 0;
        pixel_data[31][186] = 0;
        pixel_data[31][187] = 0;
        pixel_data[31][188] = 0;
        pixel_data[31][189] = 0;
        pixel_data[31][190] = 0;
        pixel_data[31][191] = 0;
        pixel_data[31][192] = 0;
        pixel_data[31][193] = 0;
        pixel_data[31][194] = 0;
        pixel_data[31][195] = 0;
        pixel_data[31][196] = 0;
        pixel_data[31][197] = 0;
        pixel_data[31][198] = 0;
        pixel_data[31][199] = 0; // y=31
        pixel_data[32][0] = 0;
        pixel_data[32][1] = 0;
        pixel_data[32][2] = 0;
        pixel_data[32][3] = 0;
        pixel_data[32][4] = 0;
        pixel_data[32][5] = 0;
        pixel_data[32][6] = 0;
        pixel_data[32][7] = 0;
        pixel_data[32][8] = 0;
        pixel_data[32][9] = 0;
        pixel_data[32][10] = 0;
        pixel_data[32][11] = 0;
        pixel_data[32][12] = 0;
        pixel_data[32][13] = 0;
        pixel_data[32][14] = 0;
        pixel_data[32][15] = 0;
        pixel_data[32][16] = 0;
        pixel_data[32][17] = 0;
        pixel_data[32][18] = 0;
        pixel_data[32][19] = 0;
        pixel_data[32][20] = 0;
        pixel_data[32][21] = 0;
        pixel_data[32][22] = 0;
        pixel_data[32][23] = 0;
        pixel_data[32][24] = 0;
        pixel_data[32][25] = 0;
        pixel_data[32][26] = 0;
        pixel_data[32][27] = 0;
        pixel_data[32][28] = 0;
        pixel_data[32][29] = 0;
        pixel_data[32][30] = 0;
        pixel_data[32][31] = 0;
        pixel_data[32][32] = 0;
        pixel_data[32][33] = 0;
        pixel_data[32][34] = 0;
        pixel_data[32][35] = 0;
        pixel_data[32][36] = 0;
        pixel_data[32][37] = 0;
        pixel_data[32][38] = 0;
        pixel_data[32][39] = 0;
        pixel_data[32][40] = 0;
        pixel_data[32][41] = 0;
        pixel_data[32][42] = 0;
        pixel_data[32][43] = 0;
        pixel_data[32][44] = 0;
        pixel_data[32][45] = 0;
        pixel_data[32][46] = 0;
        pixel_data[32][47] = 0;
        pixel_data[32][48] = 0;
        pixel_data[32][49] = 0;
        pixel_data[32][50] = 0;
        pixel_data[32][51] = 0;
        pixel_data[32][52] = 0;
        pixel_data[32][53] = 0;
        pixel_data[32][54] = 0;
        pixel_data[32][55] = 0;
        pixel_data[32][56] = 0;
        pixel_data[32][57] = 0;
        pixel_data[32][58] = 0;
        pixel_data[32][59] = 0;
        pixel_data[32][60] = 0;
        pixel_data[32][61] = 0;
        pixel_data[32][62] = 0;
        pixel_data[32][63] = 0;
        pixel_data[32][64] = 0;
        pixel_data[32][65] = 0;
        pixel_data[32][66] = 0;
        pixel_data[32][67] = 0;
        pixel_data[32][68] = 0;
        pixel_data[32][69] = 0;
        pixel_data[32][70] = 0;
        pixel_data[32][71] = 0;
        pixel_data[32][72] = 0;
        pixel_data[32][73] = 0;
        pixel_data[32][74] = 0;
        pixel_data[32][75] = 0;
        pixel_data[32][76] = 0;
        pixel_data[32][77] = 0;
        pixel_data[32][78] = 0;
        pixel_data[32][79] = 0;
        pixel_data[32][80] = 0;
        pixel_data[32][81] = 0;
        pixel_data[32][82] = 0;
        pixel_data[32][83] = 0;
        pixel_data[32][84] = 0;
        pixel_data[32][85] = 0;
        pixel_data[32][86] = 0;
        pixel_data[32][87] = 0;
        pixel_data[32][88] = 0;
        pixel_data[32][89] = 0;
        pixel_data[32][90] = 0;
        pixel_data[32][91] = 0;
        pixel_data[32][92] = 0;
        pixel_data[32][93] = 0;
        pixel_data[32][94] = 0;
        pixel_data[32][95] = 0;
        pixel_data[32][96] = 0;
        pixel_data[32][97] = 0;
        pixel_data[32][98] = 0;
        pixel_data[32][99] = 0;
        pixel_data[32][100] = 0;
        pixel_data[32][101] = 0;
        pixel_data[32][102] = 0;
        pixel_data[32][103] = 0;
        pixel_data[32][104] = 0;
        pixel_data[32][105] = 0;
        pixel_data[32][106] = 0;
        pixel_data[32][107] = 0;
        pixel_data[32][108] = 0;
        pixel_data[32][109] = 0;
        pixel_data[32][110] = 0;
        pixel_data[32][111] = 0;
        pixel_data[32][112] = 0;
        pixel_data[32][113] = 0;
        pixel_data[32][114] = 0;
        pixel_data[32][115] = 0;
        pixel_data[32][116] = 0;
        pixel_data[32][117] = 0;
        pixel_data[32][118] = 0;
        pixel_data[32][119] = 0;
        pixel_data[32][120] = 0;
        pixel_data[32][121] = 0;
        pixel_data[32][122] = 0;
        pixel_data[32][123] = 0;
        pixel_data[32][124] = 0;
        pixel_data[32][125] = 0;
        pixel_data[32][126] = 0;
        pixel_data[32][127] = 0;
        pixel_data[32][128] = 0;
        pixel_data[32][129] = 0;
        pixel_data[32][130] = 0;
        pixel_data[32][131] = 0;
        pixel_data[32][132] = 0;
        pixel_data[32][133] = 0;
        pixel_data[32][134] = 0;
        pixel_data[32][135] = 0;
        pixel_data[32][136] = 0;
        pixel_data[32][137] = 0;
        pixel_data[32][138] = 0;
        pixel_data[32][139] = 0;
        pixel_data[32][140] = 0;
        pixel_data[32][141] = 0;
        pixel_data[32][142] = 0;
        pixel_data[32][143] = 0;
        pixel_data[32][144] = 0;
        pixel_data[32][145] = 0;
        pixel_data[32][146] = 0;
        pixel_data[32][147] = 0;
        pixel_data[32][148] = 0;
        pixel_data[32][149] = 0;
        pixel_data[32][150] = 0;
        pixel_data[32][151] = 0;
        pixel_data[32][152] = 0;
        pixel_data[32][153] = 0;
        pixel_data[32][154] = 0;
        pixel_data[32][155] = 0;
        pixel_data[32][156] = 0;
        pixel_data[32][157] = 0;
        pixel_data[32][158] = 0;
        pixel_data[32][159] = 0;
        pixel_data[32][160] = 0;
        pixel_data[32][161] = 0;
        pixel_data[32][162] = 0;
        pixel_data[32][163] = 0;
        pixel_data[32][164] = 0;
        pixel_data[32][165] = 0;
        pixel_data[32][166] = 0;
        pixel_data[32][167] = 0;
        pixel_data[32][168] = 0;
        pixel_data[32][169] = 0;
        pixel_data[32][170] = 0;
        pixel_data[32][171] = 0;
        pixel_data[32][172] = 0;
        pixel_data[32][173] = 0;
        pixel_data[32][174] = 0;
        pixel_data[32][175] = 0;
        pixel_data[32][176] = 0;
        pixel_data[32][177] = 0;
        pixel_data[32][178] = 0;
        pixel_data[32][179] = 0;
        pixel_data[32][180] = 0;
        pixel_data[32][181] = 0;
        pixel_data[32][182] = 0;
        pixel_data[32][183] = 0;
        pixel_data[32][184] = 0;
        pixel_data[32][185] = 0;
        pixel_data[32][186] = 0;
        pixel_data[32][187] = 0;
        pixel_data[32][188] = 0;
        pixel_data[32][189] = 0;
        pixel_data[32][190] = 0;
        pixel_data[32][191] = 0;
        pixel_data[32][192] = 0;
        pixel_data[32][193] = 0;
        pixel_data[32][194] = 0;
        pixel_data[32][195] = 0;
        pixel_data[32][196] = 0;
        pixel_data[32][197] = 0;
        pixel_data[32][198] = 0;
        pixel_data[32][199] = 0; // y=32
        pixel_data[33][0] = 0;
        pixel_data[33][1] = 0;
        pixel_data[33][2] = 0;
        pixel_data[33][3] = 0;
        pixel_data[33][4] = 0;
        pixel_data[33][5] = 0;
        pixel_data[33][6] = 0;
        pixel_data[33][7] = 0;
        pixel_data[33][8] = 0;
        pixel_data[33][9] = 0;
        pixel_data[33][10] = 0;
        pixel_data[33][11] = 0;
        pixel_data[33][12] = 0;
        pixel_data[33][13] = 0;
        pixel_data[33][14] = 0;
        pixel_data[33][15] = 0;
        pixel_data[33][16] = 0;
        pixel_data[33][17] = 0;
        pixel_data[33][18] = 0;
        pixel_data[33][19] = 0;
        pixel_data[33][20] = 0;
        pixel_data[33][21] = 0;
        pixel_data[33][22] = 0;
        pixel_data[33][23] = 0;
        pixel_data[33][24] = 0;
        pixel_data[33][25] = 0;
        pixel_data[33][26] = 0;
        pixel_data[33][27] = 0;
        pixel_data[33][28] = 0;
        pixel_data[33][29] = 0;
        pixel_data[33][30] = 0;
        pixel_data[33][31] = 0;
        pixel_data[33][32] = 0;
        pixel_data[33][33] = 0;
        pixel_data[33][34] = 0;
        pixel_data[33][35] = 0;
        pixel_data[33][36] = 0;
        pixel_data[33][37] = 0;
        pixel_data[33][38] = 0;
        pixel_data[33][39] = 0;
        pixel_data[33][40] = 0;
        pixel_data[33][41] = 0;
        pixel_data[33][42] = 0;
        pixel_data[33][43] = 0;
        pixel_data[33][44] = 0;
        pixel_data[33][45] = 0;
        pixel_data[33][46] = 0;
        pixel_data[33][47] = 0;
        pixel_data[33][48] = 0;
        pixel_data[33][49] = 0;
        pixel_data[33][50] = 0;
        pixel_data[33][51] = 0;
        pixel_data[33][52] = 0;
        pixel_data[33][53] = 0;
        pixel_data[33][54] = 0;
        pixel_data[33][55] = 0;
        pixel_data[33][56] = 0;
        pixel_data[33][57] = 0;
        pixel_data[33][58] = 0;
        pixel_data[33][59] = 0;
        pixel_data[33][60] = 0;
        pixel_data[33][61] = 0;
        pixel_data[33][62] = 0;
        pixel_data[33][63] = 0;
        pixel_data[33][64] = 0;
        pixel_data[33][65] = 0;
        pixel_data[33][66] = 0;
        pixel_data[33][67] = 0;
        pixel_data[33][68] = 0;
        pixel_data[33][69] = 0;
        pixel_data[33][70] = 0;
        pixel_data[33][71] = 0;
        pixel_data[33][72] = 0;
        pixel_data[33][73] = 0;
        pixel_data[33][74] = 0;
        pixel_data[33][75] = 0;
        pixel_data[33][76] = 0;
        pixel_data[33][77] = 0;
        pixel_data[33][78] = 0;
        pixel_data[33][79] = 0;
        pixel_data[33][80] = 0;
        pixel_data[33][81] = 0;
        pixel_data[33][82] = 0;
        pixel_data[33][83] = 0;
        pixel_data[33][84] = 0;
        pixel_data[33][85] = 0;
        pixel_data[33][86] = 0;
        pixel_data[33][87] = 0;
        pixel_data[33][88] = 0;
        pixel_data[33][89] = 0;
        pixel_data[33][90] = 0;
        pixel_data[33][91] = 0;
        pixel_data[33][92] = 0;
        pixel_data[33][93] = 0;
        pixel_data[33][94] = 0;
        pixel_data[33][95] = 0;
        pixel_data[33][96] = 0;
        pixel_data[33][97] = 0;
        pixel_data[33][98] = 0;
        pixel_data[33][99] = 0;
        pixel_data[33][100] = 0;
        pixel_data[33][101] = 0;
        pixel_data[33][102] = 0;
        pixel_data[33][103] = 0;
        pixel_data[33][104] = 0;
        pixel_data[33][105] = 0;
        pixel_data[33][106] = 0;
        pixel_data[33][107] = 0;
        pixel_data[33][108] = 0;
        pixel_data[33][109] = 0;
        pixel_data[33][110] = 0;
        pixel_data[33][111] = 0;
        pixel_data[33][112] = 0;
        pixel_data[33][113] = 0;
        pixel_data[33][114] = 0;
        pixel_data[33][115] = 0;
        pixel_data[33][116] = 0;
        pixel_data[33][117] = 0;
        pixel_data[33][118] = 0;
        pixel_data[33][119] = 0;
        pixel_data[33][120] = 0;
        pixel_data[33][121] = 0;
        pixel_data[33][122] = 0;
        pixel_data[33][123] = 0;
        pixel_data[33][124] = 0;
        pixel_data[33][125] = 0;
        pixel_data[33][126] = 0;
        pixel_data[33][127] = 0;
        pixel_data[33][128] = 0;
        pixel_data[33][129] = 0;
        pixel_data[33][130] = 0;
        pixel_data[33][131] = 0;
        pixel_data[33][132] = 0;
        pixel_data[33][133] = 0;
        pixel_data[33][134] = 0;
        pixel_data[33][135] = 0;
        pixel_data[33][136] = 0;
        pixel_data[33][137] = 0;
        pixel_data[33][138] = 0;
        pixel_data[33][139] = 0;
        pixel_data[33][140] = 0;
        pixel_data[33][141] = 0;
        pixel_data[33][142] = 0;
        pixel_data[33][143] = 0;
        pixel_data[33][144] = 0;
        pixel_data[33][145] = 0;
        pixel_data[33][146] = 0;
        pixel_data[33][147] = 0;
        pixel_data[33][148] = 0;
        pixel_data[33][149] = 0;
        pixel_data[33][150] = 0;
        pixel_data[33][151] = 0;
        pixel_data[33][152] = 0;
        pixel_data[33][153] = 0;
        pixel_data[33][154] = 0;
        pixel_data[33][155] = 0;
        pixel_data[33][156] = 0;
        pixel_data[33][157] = 0;
        pixel_data[33][158] = 0;
        pixel_data[33][159] = 0;
        pixel_data[33][160] = 0;
        pixel_data[33][161] = 0;
        pixel_data[33][162] = 0;
        pixel_data[33][163] = 0;
        pixel_data[33][164] = 0;
        pixel_data[33][165] = 0;
        pixel_data[33][166] = 0;
        pixel_data[33][167] = 0;
        pixel_data[33][168] = 0;
        pixel_data[33][169] = 0;
        pixel_data[33][170] = 0;
        pixel_data[33][171] = 0;
        pixel_data[33][172] = 0;
        pixel_data[33][173] = 0;
        pixel_data[33][174] = 0;
        pixel_data[33][175] = 0;
        pixel_data[33][176] = 0;
        pixel_data[33][177] = 0;
        pixel_data[33][178] = 0;
        pixel_data[33][179] = 0;
        pixel_data[33][180] = 0;
        pixel_data[33][181] = 0;
        pixel_data[33][182] = 0;
        pixel_data[33][183] = 0;
        pixel_data[33][184] = 0;
        pixel_data[33][185] = 0;
        pixel_data[33][186] = 0;
        pixel_data[33][187] = 0;
        pixel_data[33][188] = 0;
        pixel_data[33][189] = 0;
        pixel_data[33][190] = 0;
        pixel_data[33][191] = 0;
        pixel_data[33][192] = 0;
        pixel_data[33][193] = 0;
        pixel_data[33][194] = 0;
        pixel_data[33][195] = 0;
        pixel_data[33][196] = 0;
        pixel_data[33][197] = 0;
        pixel_data[33][198] = 0;
        pixel_data[33][199] = 0; // y=33
        pixel_data[34][0] = 0;
        pixel_data[34][1] = 0;
        pixel_data[34][2] = 0;
        pixel_data[34][3] = 0;
        pixel_data[34][4] = 0;
        pixel_data[34][5] = 0;
        pixel_data[34][6] = 0;
        pixel_data[34][7] = 0;
        pixel_data[34][8] = 0;
        pixel_data[34][9] = 0;
        pixel_data[34][10] = 0;
        pixel_data[34][11] = 0;
        pixel_data[34][12] = 0;
        pixel_data[34][13] = 0;
        pixel_data[34][14] = 0;
        pixel_data[34][15] = 0;
        pixel_data[34][16] = 0;
        pixel_data[34][17] = 0;
        pixel_data[34][18] = 0;
        pixel_data[34][19] = 0;
        pixel_data[34][20] = 0;
        pixel_data[34][21] = 0;
        pixel_data[34][22] = 0;
        pixel_data[34][23] = 0;
        pixel_data[34][24] = 0;
        pixel_data[34][25] = 0;
        pixel_data[34][26] = 0;
        pixel_data[34][27] = 0;
        pixel_data[34][28] = 0;
        pixel_data[34][29] = 0;
        pixel_data[34][30] = 0;
        pixel_data[34][31] = 0;
        pixel_data[34][32] = 0;
        pixel_data[34][33] = 0;
        pixel_data[34][34] = 0;
        pixel_data[34][35] = 0;
        pixel_data[34][36] = 0;
        pixel_data[34][37] = 0;
        pixel_data[34][38] = 0;
        pixel_data[34][39] = 0;
        pixel_data[34][40] = 0;
        pixel_data[34][41] = 0;
        pixel_data[34][42] = 0;
        pixel_data[34][43] = 0;
        pixel_data[34][44] = 0;
        pixel_data[34][45] = 0;
        pixel_data[34][46] = 0;
        pixel_data[34][47] = 0;
        pixel_data[34][48] = 0;
        pixel_data[34][49] = 0;
        pixel_data[34][50] = 0;
        pixel_data[34][51] = 0;
        pixel_data[34][52] = 0;
        pixel_data[34][53] = 0;
        pixel_data[34][54] = 0;
        pixel_data[34][55] = 0;
        pixel_data[34][56] = 0;
        pixel_data[34][57] = 0;
        pixel_data[34][58] = 0;
        pixel_data[34][59] = 0;
        pixel_data[34][60] = 0;
        pixel_data[34][61] = 0;
        pixel_data[34][62] = 0;
        pixel_data[34][63] = 0;
        pixel_data[34][64] = 0;
        pixel_data[34][65] = 0;
        pixel_data[34][66] = 0;
        pixel_data[34][67] = 0;
        pixel_data[34][68] = 0;
        pixel_data[34][69] = 0;
        pixel_data[34][70] = 0;
        pixel_data[34][71] = 0;
        pixel_data[34][72] = 0;
        pixel_data[34][73] = 0;
        pixel_data[34][74] = 0;
        pixel_data[34][75] = 0;
        pixel_data[34][76] = 0;
        pixel_data[34][77] = 0;
        pixel_data[34][78] = 0;
        pixel_data[34][79] = 0;
        pixel_data[34][80] = 0;
        pixel_data[34][81] = 0;
        pixel_data[34][82] = 0;
        pixel_data[34][83] = 0;
        pixel_data[34][84] = 0;
        pixel_data[34][85] = 0;
        pixel_data[34][86] = 0;
        pixel_data[34][87] = 0;
        pixel_data[34][88] = 0;
        pixel_data[34][89] = 0;
        pixel_data[34][90] = 0;
        pixel_data[34][91] = 0;
        pixel_data[34][92] = 0;
        pixel_data[34][93] = 0;
        pixel_data[34][94] = 0;
        pixel_data[34][95] = 0;
        pixel_data[34][96] = 0;
        pixel_data[34][97] = 0;
        pixel_data[34][98] = 0;
        pixel_data[34][99] = 0;
        pixel_data[34][100] = 0;
        pixel_data[34][101] = 0;
        pixel_data[34][102] = 0;
        pixel_data[34][103] = 0;
        pixel_data[34][104] = 0;
        pixel_data[34][105] = 0;
        pixel_data[34][106] = 0;
        pixel_data[34][107] = 0;
        pixel_data[34][108] = 0;
        pixel_data[34][109] = 0;
        pixel_data[34][110] = 0;
        pixel_data[34][111] = 0;
        pixel_data[34][112] = 0;
        pixel_data[34][113] = 0;
        pixel_data[34][114] = 0;
        pixel_data[34][115] = 0;
        pixel_data[34][116] = 0;
        pixel_data[34][117] = 0;
        pixel_data[34][118] = 0;
        pixel_data[34][119] = 0;
        pixel_data[34][120] = 0;
        pixel_data[34][121] = 0;
        pixel_data[34][122] = 0;
        pixel_data[34][123] = 0;
        pixel_data[34][124] = 0;
        pixel_data[34][125] = 0;
        pixel_data[34][126] = 0;
        pixel_data[34][127] = 0;
        pixel_data[34][128] = 0;
        pixel_data[34][129] = 0;
        pixel_data[34][130] = 0;
        pixel_data[34][131] = 0;
        pixel_data[34][132] = 0;
        pixel_data[34][133] = 0;
        pixel_data[34][134] = 0;
        pixel_data[34][135] = 0;
        pixel_data[34][136] = 0;
        pixel_data[34][137] = 0;
        pixel_data[34][138] = 0;
        pixel_data[34][139] = 0;
        pixel_data[34][140] = 0;
        pixel_data[34][141] = 0;
        pixel_data[34][142] = 0;
        pixel_data[34][143] = 0;
        pixel_data[34][144] = 0;
        pixel_data[34][145] = 0;
        pixel_data[34][146] = 0;
        pixel_data[34][147] = 0;
        pixel_data[34][148] = 0;
        pixel_data[34][149] = 0;
        pixel_data[34][150] = 0;
        pixel_data[34][151] = 0;
        pixel_data[34][152] = 0;
        pixel_data[34][153] = 0;
        pixel_data[34][154] = 0;
        pixel_data[34][155] = 0;
        pixel_data[34][156] = 0;
        pixel_data[34][157] = 0;
        pixel_data[34][158] = 0;
        pixel_data[34][159] = 0;
        pixel_data[34][160] = 0;
        pixel_data[34][161] = 0;
        pixel_data[34][162] = 0;
        pixel_data[34][163] = 0;
        pixel_data[34][164] = 0;
        pixel_data[34][165] = 0;
        pixel_data[34][166] = 0;
        pixel_data[34][167] = 0;
        pixel_data[34][168] = 0;
        pixel_data[34][169] = 0;
        pixel_data[34][170] = 0;
        pixel_data[34][171] = 0;
        pixel_data[34][172] = 0;
        pixel_data[34][173] = 0;
        pixel_data[34][174] = 0;
        pixel_data[34][175] = 0;
        pixel_data[34][176] = 0;
        pixel_data[34][177] = 0;
        pixel_data[34][178] = 0;
        pixel_data[34][179] = 0;
        pixel_data[34][180] = 0;
        pixel_data[34][181] = 0;
        pixel_data[34][182] = 0;
        pixel_data[34][183] = 0;
        pixel_data[34][184] = 0;
        pixel_data[34][185] = 0;
        pixel_data[34][186] = 0;
        pixel_data[34][187] = 0;
        pixel_data[34][188] = 0;
        pixel_data[34][189] = 0;
        pixel_data[34][190] = 0;
        pixel_data[34][191] = 0;
        pixel_data[34][192] = 0;
        pixel_data[34][193] = 0;
        pixel_data[34][194] = 0;
        pixel_data[34][195] = 0;
        pixel_data[34][196] = 0;
        pixel_data[34][197] = 0;
        pixel_data[34][198] = 0;
        pixel_data[34][199] = 0; // y=34
        pixel_data[35][0] = 0;
        pixel_data[35][1] = 0;
        pixel_data[35][2] = 0;
        pixel_data[35][3] = 0;
        pixel_data[35][4] = 0;
        pixel_data[35][5] = 0;
        pixel_data[35][6] = 0;
        pixel_data[35][7] = 0;
        pixel_data[35][8] = 0;
        pixel_data[35][9] = 0;
        pixel_data[35][10] = 0;
        pixel_data[35][11] = 0;
        pixel_data[35][12] = 0;
        pixel_data[35][13] = 0;
        pixel_data[35][14] = 0;
        pixel_data[35][15] = 0;
        pixel_data[35][16] = 0;
        pixel_data[35][17] = 0;
        pixel_data[35][18] = 0;
        pixel_data[35][19] = 0;
        pixel_data[35][20] = 0;
        pixel_data[35][21] = 0;
        pixel_data[35][22] = 0;
        pixel_data[35][23] = 0;
        pixel_data[35][24] = 0;
        pixel_data[35][25] = 0;
        pixel_data[35][26] = 0;
        pixel_data[35][27] = 0;
        pixel_data[35][28] = 0;
        pixel_data[35][29] = 0;
        pixel_data[35][30] = 0;
        pixel_data[35][31] = 0;
        pixel_data[35][32] = 0;
        pixel_data[35][33] = 0;
        pixel_data[35][34] = 0;
        pixel_data[35][35] = 0;
        pixel_data[35][36] = 0;
        pixel_data[35][37] = 0;
        pixel_data[35][38] = 0;
        pixel_data[35][39] = 0;
        pixel_data[35][40] = 0;
        pixel_data[35][41] = 0;
        pixel_data[35][42] = 0;
        pixel_data[35][43] = 0;
        pixel_data[35][44] = 0;
        pixel_data[35][45] = 0;
        pixel_data[35][46] = 0;
        pixel_data[35][47] = 0;
        pixel_data[35][48] = 0;
        pixel_data[35][49] = 0;
        pixel_data[35][50] = 0;
        pixel_data[35][51] = 0;
        pixel_data[35][52] = 0;
        pixel_data[35][53] = 0;
        pixel_data[35][54] = 0;
        pixel_data[35][55] = 0;
        pixel_data[35][56] = 0;
        pixel_data[35][57] = 0;
        pixel_data[35][58] = 0;
        pixel_data[35][59] = 0;
        pixel_data[35][60] = 0;
        pixel_data[35][61] = 0;
        pixel_data[35][62] = 0;
        pixel_data[35][63] = 0;
        pixel_data[35][64] = 0;
        pixel_data[35][65] = 0;
        pixel_data[35][66] = 0;
        pixel_data[35][67] = 0;
        pixel_data[35][68] = 0;
        pixel_data[35][69] = 0;
        pixel_data[35][70] = 0;
        pixel_data[35][71] = 0;
        pixel_data[35][72] = 0;
        pixel_data[35][73] = 0;
        pixel_data[35][74] = 0;
        pixel_data[35][75] = 0;
        pixel_data[35][76] = 0;
        pixel_data[35][77] = 0;
        pixel_data[35][78] = 0;
        pixel_data[35][79] = 0;
        pixel_data[35][80] = 0;
        pixel_data[35][81] = 0;
        pixel_data[35][82] = 0;
        pixel_data[35][83] = 0;
        pixel_data[35][84] = 0;
        pixel_data[35][85] = 0;
        pixel_data[35][86] = 0;
        pixel_data[35][87] = 0;
        pixel_data[35][88] = 0;
        pixel_data[35][89] = 0;
        pixel_data[35][90] = 0;
        pixel_data[35][91] = 0;
        pixel_data[35][92] = 0;
        pixel_data[35][93] = 0;
        pixel_data[35][94] = 0;
        pixel_data[35][95] = 0;
        pixel_data[35][96] = 0;
        pixel_data[35][97] = 0;
        pixel_data[35][98] = 0;
        pixel_data[35][99] = 0;
        pixel_data[35][100] = 0;
        pixel_data[35][101] = 0;
        pixel_data[35][102] = 0;
        pixel_data[35][103] = 0;
        pixel_data[35][104] = 0;
        pixel_data[35][105] = 0;
        pixel_data[35][106] = 0;
        pixel_data[35][107] = 0;
        pixel_data[35][108] = 0;
        pixel_data[35][109] = 0;
        pixel_data[35][110] = 0;
        pixel_data[35][111] = 0;
        pixel_data[35][112] = 0;
        pixel_data[35][113] = 0;
        pixel_data[35][114] = 0;
        pixel_data[35][115] = 0;
        pixel_data[35][116] = 0;
        pixel_data[35][117] = 0;
        pixel_data[35][118] = 0;
        pixel_data[35][119] = 0;
        pixel_data[35][120] = 0;
        pixel_data[35][121] = 0;
        pixel_data[35][122] = 0;
        pixel_data[35][123] = 0;
        pixel_data[35][124] = 0;
        pixel_data[35][125] = 0;
        pixel_data[35][126] = 0;
        pixel_data[35][127] = 0;
        pixel_data[35][128] = 0;
        pixel_data[35][129] = 0;
        pixel_data[35][130] = 0;
        pixel_data[35][131] = 0;
        pixel_data[35][132] = 0;
        pixel_data[35][133] = 0;
        pixel_data[35][134] = 0;
        pixel_data[35][135] = 0;
        pixel_data[35][136] = 0;
        pixel_data[35][137] = 0;
        pixel_data[35][138] = 0;
        pixel_data[35][139] = 0;
        pixel_data[35][140] = 0;
        pixel_data[35][141] = 0;
        pixel_data[35][142] = 0;
        pixel_data[35][143] = 0;
        pixel_data[35][144] = 0;
        pixel_data[35][145] = 0;
        pixel_data[35][146] = 0;
        pixel_data[35][147] = 0;
        pixel_data[35][148] = 0;
        pixel_data[35][149] = 0;
        pixel_data[35][150] = 0;
        pixel_data[35][151] = 0;
        pixel_data[35][152] = 0;
        pixel_data[35][153] = 0;
        pixel_data[35][154] = 0;
        pixel_data[35][155] = 0;
        pixel_data[35][156] = 0;
        pixel_data[35][157] = 0;
        pixel_data[35][158] = 0;
        pixel_data[35][159] = 0;
        pixel_data[35][160] = 0;
        pixel_data[35][161] = 0;
        pixel_data[35][162] = 0;
        pixel_data[35][163] = 0;
        pixel_data[35][164] = 0;
        pixel_data[35][165] = 0;
        pixel_data[35][166] = 0;
        pixel_data[35][167] = 0;
        pixel_data[35][168] = 0;
        pixel_data[35][169] = 0;
        pixel_data[35][170] = 0;
        pixel_data[35][171] = 0;
        pixel_data[35][172] = 0;
        pixel_data[35][173] = 0;
        pixel_data[35][174] = 0;
        pixel_data[35][175] = 0;
        pixel_data[35][176] = 0;
        pixel_data[35][177] = 0;
        pixel_data[35][178] = 0;
        pixel_data[35][179] = 0;
        pixel_data[35][180] = 0;
        pixel_data[35][181] = 0;
        pixel_data[35][182] = 0;
        pixel_data[35][183] = 0;
        pixel_data[35][184] = 0;
        pixel_data[35][185] = 0;
        pixel_data[35][186] = 0;
        pixel_data[35][187] = 0;
        pixel_data[35][188] = 0;
        pixel_data[35][189] = 0;
        pixel_data[35][190] = 0;
        pixel_data[35][191] = 0;
        pixel_data[35][192] = 0;
        pixel_data[35][193] = 0;
        pixel_data[35][194] = 0;
        pixel_data[35][195] = 0;
        pixel_data[35][196] = 0;
        pixel_data[35][197] = 0;
        pixel_data[35][198] = 0;
        pixel_data[35][199] = 0; // y=35
        pixel_data[36][0] = 0;
        pixel_data[36][1] = 0;
        pixel_data[36][2] = 0;
        pixel_data[36][3] = 0;
        pixel_data[36][4] = 0;
        pixel_data[36][5] = 0;
        pixel_data[36][6] = 0;
        pixel_data[36][7] = 0;
        pixel_data[36][8] = 0;
        pixel_data[36][9] = 0;
        pixel_data[36][10] = 0;
        pixel_data[36][11] = 0;
        pixel_data[36][12] = 0;
        pixel_data[36][13] = 0;
        pixel_data[36][14] = 0;
        pixel_data[36][15] = 0;
        pixel_data[36][16] = 0;
        pixel_data[36][17] = 0;
        pixel_data[36][18] = 0;
        pixel_data[36][19] = 0;
        pixel_data[36][20] = 0;
        pixel_data[36][21] = 0;
        pixel_data[36][22] = 0;
        pixel_data[36][23] = 0;
        pixel_data[36][24] = 0;
        pixel_data[36][25] = 0;
        pixel_data[36][26] = 0;
        pixel_data[36][27] = 0;
        pixel_data[36][28] = 0;
        pixel_data[36][29] = 0;
        pixel_data[36][30] = 0;
        pixel_data[36][31] = 0;
        pixel_data[36][32] = 0;
        pixel_data[36][33] = 0;
        pixel_data[36][34] = 0;
        pixel_data[36][35] = 0;
        pixel_data[36][36] = 0;
        pixel_data[36][37] = 0;
        pixel_data[36][38] = 0;
        pixel_data[36][39] = 0;
        pixel_data[36][40] = 0;
        pixel_data[36][41] = 0;
        pixel_data[36][42] = 0;
        pixel_data[36][43] = 0;
        pixel_data[36][44] = 0;
        pixel_data[36][45] = 0;
        pixel_data[36][46] = 0;
        pixel_data[36][47] = 0;
        pixel_data[36][48] = 0;
        pixel_data[36][49] = 0;
        pixel_data[36][50] = 0;
        pixel_data[36][51] = 0;
        pixel_data[36][52] = 0;
        pixel_data[36][53] = 0;
        pixel_data[36][54] = 0;
        pixel_data[36][55] = 0;
        pixel_data[36][56] = 0;
        pixel_data[36][57] = 0;
        pixel_data[36][58] = 0;
        pixel_data[36][59] = 0;
        pixel_data[36][60] = 0;
        pixel_data[36][61] = 0;
        pixel_data[36][62] = 0;
        pixel_data[36][63] = 0;
        pixel_data[36][64] = 0;
        pixel_data[36][65] = 0;
        pixel_data[36][66] = 0;
        pixel_data[36][67] = 0;
        pixel_data[36][68] = 0;
        pixel_data[36][69] = 0;
        pixel_data[36][70] = 0;
        pixel_data[36][71] = 0;
        pixel_data[36][72] = 0;
        pixel_data[36][73] = 0;
        pixel_data[36][74] = 0;
        pixel_data[36][75] = 0;
        pixel_data[36][76] = 0;
        pixel_data[36][77] = 0;
        pixel_data[36][78] = 0;
        pixel_data[36][79] = 0;
        pixel_data[36][80] = 0;
        pixel_data[36][81] = 0;
        pixel_data[36][82] = 0;
        pixel_data[36][83] = 0;
        pixel_data[36][84] = 0;
        pixel_data[36][85] = 0;
        pixel_data[36][86] = 0;
        pixel_data[36][87] = 0;
        pixel_data[36][88] = 0;
        pixel_data[36][89] = 0;
        pixel_data[36][90] = 0;
        pixel_data[36][91] = 0;
        pixel_data[36][92] = 0;
        pixel_data[36][93] = 0;
        pixel_data[36][94] = 0;
        pixel_data[36][95] = 0;
        pixel_data[36][96] = 0;
        pixel_data[36][97] = 0;
        pixel_data[36][98] = 0;
        pixel_data[36][99] = 0;
        pixel_data[36][100] = 0;
        pixel_data[36][101] = 0;
        pixel_data[36][102] = 0;
        pixel_data[36][103] = 0;
        pixel_data[36][104] = 0;
        pixel_data[36][105] = 0;
        pixel_data[36][106] = 0;
        pixel_data[36][107] = 0;
        pixel_data[36][108] = 0;
        pixel_data[36][109] = 0;
        pixel_data[36][110] = 0;
        pixel_data[36][111] = 0;
        pixel_data[36][112] = 0;
        pixel_data[36][113] = 0;
        pixel_data[36][114] = 0;
        pixel_data[36][115] = 0;
        pixel_data[36][116] = 0;
        pixel_data[36][117] = 0;
        pixel_data[36][118] = 0;
        pixel_data[36][119] = 0;
        pixel_data[36][120] = 0;
        pixel_data[36][121] = 0;
        pixel_data[36][122] = 0;
        pixel_data[36][123] = 0;
        pixel_data[36][124] = 0;
        pixel_data[36][125] = 0;
        pixel_data[36][126] = 0;
        pixel_data[36][127] = 0;
        pixel_data[36][128] = 0;
        pixel_data[36][129] = 0;
        pixel_data[36][130] = 0;
        pixel_data[36][131] = 0;
        pixel_data[36][132] = 0;
        pixel_data[36][133] = 0;
        pixel_data[36][134] = 0;
        pixel_data[36][135] = 0;
        pixel_data[36][136] = 0;
        pixel_data[36][137] = 0;
        pixel_data[36][138] = 0;
        pixel_data[36][139] = 0;
        pixel_data[36][140] = 0;
        pixel_data[36][141] = 0;
        pixel_data[36][142] = 0;
        pixel_data[36][143] = 0;
        pixel_data[36][144] = 0;
        pixel_data[36][145] = 0;
        pixel_data[36][146] = 0;
        pixel_data[36][147] = 0;
        pixel_data[36][148] = 0;
        pixel_data[36][149] = 0;
        pixel_data[36][150] = 0;
        pixel_data[36][151] = 0;
        pixel_data[36][152] = 0;
        pixel_data[36][153] = 0;
        pixel_data[36][154] = 0;
        pixel_data[36][155] = 0;
        pixel_data[36][156] = 0;
        pixel_data[36][157] = 0;
        pixel_data[36][158] = 0;
        pixel_data[36][159] = 0;
        pixel_data[36][160] = 0;
        pixel_data[36][161] = 0;
        pixel_data[36][162] = 0;
        pixel_data[36][163] = 0;
        pixel_data[36][164] = 0;
        pixel_data[36][165] = 0;
        pixel_data[36][166] = 0;
        pixel_data[36][167] = 0;
        pixel_data[36][168] = 0;
        pixel_data[36][169] = 0;
        pixel_data[36][170] = 0;
        pixel_data[36][171] = 0;
        pixel_data[36][172] = 0;
        pixel_data[36][173] = 0;
        pixel_data[36][174] = 0;
        pixel_data[36][175] = 0;
        pixel_data[36][176] = 0;
        pixel_data[36][177] = 0;
        pixel_data[36][178] = 0;
        pixel_data[36][179] = 0;
        pixel_data[36][180] = 0;
        pixel_data[36][181] = 0;
        pixel_data[36][182] = 0;
        pixel_data[36][183] = 0;
        pixel_data[36][184] = 0;
        pixel_data[36][185] = 0;
        pixel_data[36][186] = 0;
        pixel_data[36][187] = 0;
        pixel_data[36][188] = 0;
        pixel_data[36][189] = 0;
        pixel_data[36][190] = 0;
        pixel_data[36][191] = 0;
        pixel_data[36][192] = 0;
        pixel_data[36][193] = 0;
        pixel_data[36][194] = 0;
        pixel_data[36][195] = 0;
        pixel_data[36][196] = 0;
        pixel_data[36][197] = 0;
        pixel_data[36][198] = 0;
        pixel_data[36][199] = 0; // y=36
        pixel_data[37][0] = 0;
        pixel_data[37][1] = 0;
        pixel_data[37][2] = 0;
        pixel_data[37][3] = 0;
        pixel_data[37][4] = 0;
        pixel_data[37][5] = 0;
        pixel_data[37][6] = 0;
        pixel_data[37][7] = 0;
        pixel_data[37][8] = 0;
        pixel_data[37][9] = 0;
        pixel_data[37][10] = 0;
        pixel_data[37][11] = 0;
        pixel_data[37][12] = 0;
        pixel_data[37][13] = 0;
        pixel_data[37][14] = 0;
        pixel_data[37][15] = 0;
        pixel_data[37][16] = 0;
        pixel_data[37][17] = 0;
        pixel_data[37][18] = 0;
        pixel_data[37][19] = 0;
        pixel_data[37][20] = 0;
        pixel_data[37][21] = 0;
        pixel_data[37][22] = 0;
        pixel_data[37][23] = 0;
        pixel_data[37][24] = 0;
        pixel_data[37][25] = 0;
        pixel_data[37][26] = 0;
        pixel_data[37][27] = 0;
        pixel_data[37][28] = 0;
        pixel_data[37][29] = 0;
        pixel_data[37][30] = 0;
        pixel_data[37][31] = 0;
        pixel_data[37][32] = 0;
        pixel_data[37][33] = 0;
        pixel_data[37][34] = 0;
        pixel_data[37][35] = 0;
        pixel_data[37][36] = 0;
        pixel_data[37][37] = 0;
        pixel_data[37][38] = 0;
        pixel_data[37][39] = 0;
        pixel_data[37][40] = 0;
        pixel_data[37][41] = 0;
        pixel_data[37][42] = 0;
        pixel_data[37][43] = 0;
        pixel_data[37][44] = 0;
        pixel_data[37][45] = 0;
        pixel_data[37][46] = 0;
        pixel_data[37][47] = 0;
        pixel_data[37][48] = 0;
        pixel_data[37][49] = 0;
        pixel_data[37][50] = 0;
        pixel_data[37][51] = 0;
        pixel_data[37][52] = 0;
        pixel_data[37][53] = 0;
        pixel_data[37][54] = 0;
        pixel_data[37][55] = 0;
        pixel_data[37][56] = 0;
        pixel_data[37][57] = 0;
        pixel_data[37][58] = 0;
        pixel_data[37][59] = 0;
        pixel_data[37][60] = 0;
        pixel_data[37][61] = 0;
        pixel_data[37][62] = 0;
        pixel_data[37][63] = 0;
        pixel_data[37][64] = 0;
        pixel_data[37][65] = 0;
        pixel_data[37][66] = 0;
        pixel_data[37][67] = 0;
        pixel_data[37][68] = 0;
        pixel_data[37][69] = 0;
        pixel_data[37][70] = 0;
        pixel_data[37][71] = 0;
        pixel_data[37][72] = 0;
        pixel_data[37][73] = 0;
        pixel_data[37][74] = 0;
        pixel_data[37][75] = 0;
        pixel_data[37][76] = 0;
        pixel_data[37][77] = 0;
        pixel_data[37][78] = 0;
        pixel_data[37][79] = 0;
        pixel_data[37][80] = 0;
        pixel_data[37][81] = 0;
        pixel_data[37][82] = 0;
        pixel_data[37][83] = 0;
        pixel_data[37][84] = 0;
        pixel_data[37][85] = 0;
        pixel_data[37][86] = 0;
        pixel_data[37][87] = 0;
        pixel_data[37][88] = 0;
        pixel_data[37][89] = 0;
        pixel_data[37][90] = 0;
        pixel_data[37][91] = 0;
        pixel_data[37][92] = 0;
        pixel_data[37][93] = 0;
        pixel_data[37][94] = 0;
        pixel_data[37][95] = 0;
        pixel_data[37][96] = 0;
        pixel_data[37][97] = 0;
        pixel_data[37][98] = 0;
        pixel_data[37][99] = 0;
        pixel_data[37][100] = 0;
        pixel_data[37][101] = 0;
        pixel_data[37][102] = 0;
        pixel_data[37][103] = 0;
        pixel_data[37][104] = 0;
        pixel_data[37][105] = 0;
        pixel_data[37][106] = 0;
        pixel_data[37][107] = 0;
        pixel_data[37][108] = 0;
        pixel_data[37][109] = 0;
        pixel_data[37][110] = 0;
        pixel_data[37][111] = 0;
        pixel_data[37][112] = 0;
        pixel_data[37][113] = 0;
        pixel_data[37][114] = 0;
        pixel_data[37][115] = 0;
        pixel_data[37][116] = 0;
        pixel_data[37][117] = 0;
        pixel_data[37][118] = 0;
        pixel_data[37][119] = 0;
        pixel_data[37][120] = 0;
        pixel_data[37][121] = 0;
        pixel_data[37][122] = 0;
        pixel_data[37][123] = 0;
        pixel_data[37][124] = 0;
        pixel_data[37][125] = 0;
        pixel_data[37][126] = 0;
        pixel_data[37][127] = 0;
        pixel_data[37][128] = 0;
        pixel_data[37][129] = 0;
        pixel_data[37][130] = 0;
        pixel_data[37][131] = 0;
        pixel_data[37][132] = 0;
        pixel_data[37][133] = 0;
        pixel_data[37][134] = 0;
        pixel_data[37][135] = 0;
        pixel_data[37][136] = 0;
        pixel_data[37][137] = 0;
        pixel_data[37][138] = 0;
        pixel_data[37][139] = 0;
        pixel_data[37][140] = 0;
        pixel_data[37][141] = 0;
        pixel_data[37][142] = 0;
        pixel_data[37][143] = 0;
        pixel_data[37][144] = 0;
        pixel_data[37][145] = 0;
        pixel_data[37][146] = 0;
        pixel_data[37][147] = 0;
        pixel_data[37][148] = 0;
        pixel_data[37][149] = 0;
        pixel_data[37][150] = 0;
        pixel_data[37][151] = 0;
        pixel_data[37][152] = 0;
        pixel_data[37][153] = 0;
        pixel_data[37][154] = 0;
        pixel_data[37][155] = 0;
        pixel_data[37][156] = 0;
        pixel_data[37][157] = 0;
        pixel_data[37][158] = 0;
        pixel_data[37][159] = 0;
        pixel_data[37][160] = 0;
        pixel_data[37][161] = 0;
        pixel_data[37][162] = 0;
        pixel_data[37][163] = 0;
        pixel_data[37][164] = 0;
        pixel_data[37][165] = 0;
        pixel_data[37][166] = 0;
        pixel_data[37][167] = 0;
        pixel_data[37][168] = 0;
        pixel_data[37][169] = 0;
        pixel_data[37][170] = 0;
        pixel_data[37][171] = 0;
        pixel_data[37][172] = 0;
        pixel_data[37][173] = 0;
        pixel_data[37][174] = 0;
        pixel_data[37][175] = 0;
        pixel_data[37][176] = 0;
        pixel_data[37][177] = 0;
        pixel_data[37][178] = 0;
        pixel_data[37][179] = 0;
        pixel_data[37][180] = 0;
        pixel_data[37][181] = 0;
        pixel_data[37][182] = 0;
        pixel_data[37][183] = 0;
        pixel_data[37][184] = 0;
        pixel_data[37][185] = 0;
        pixel_data[37][186] = 0;
        pixel_data[37][187] = 0;
        pixel_data[37][188] = 0;
        pixel_data[37][189] = 0;
        pixel_data[37][190] = 0;
        pixel_data[37][191] = 0;
        pixel_data[37][192] = 0;
        pixel_data[37][193] = 0;
        pixel_data[37][194] = 0;
        pixel_data[37][195] = 0;
        pixel_data[37][196] = 0;
        pixel_data[37][197] = 0;
        pixel_data[37][198] = 0;
        pixel_data[37][199] = 0; // y=37
        pixel_data[38][0] = 0;
        pixel_data[38][1] = 0;
        pixel_data[38][2] = 0;
        pixel_data[38][3] = 0;
        pixel_data[38][4] = 0;
        pixel_data[38][5] = 0;
        pixel_data[38][6] = 0;
        pixel_data[38][7] = 0;
        pixel_data[38][8] = 0;
        pixel_data[38][9] = 0;
        pixel_data[38][10] = 0;
        pixel_data[38][11] = 0;
        pixel_data[38][12] = 0;
        pixel_data[38][13] = 0;
        pixel_data[38][14] = 0;
        pixel_data[38][15] = 0;
        pixel_data[38][16] = 0;
        pixel_data[38][17] = 0;
        pixel_data[38][18] = 0;
        pixel_data[38][19] = 0;
        pixel_data[38][20] = 0;
        pixel_data[38][21] = 0;
        pixel_data[38][22] = 0;
        pixel_data[38][23] = 0;
        pixel_data[38][24] = 0;
        pixel_data[38][25] = 0;
        pixel_data[38][26] = 0;
        pixel_data[38][27] = 0;
        pixel_data[38][28] = 0;
        pixel_data[38][29] = 0;
        pixel_data[38][30] = 0;
        pixel_data[38][31] = 0;
        pixel_data[38][32] = 0;
        pixel_data[38][33] = 0;
        pixel_data[38][34] = 0;
        pixel_data[38][35] = 0;
        pixel_data[38][36] = 0;
        pixel_data[38][37] = 0;
        pixel_data[38][38] = 0;
        pixel_data[38][39] = 0;
        pixel_data[38][40] = 0;
        pixel_data[38][41] = 0;
        pixel_data[38][42] = 0;
        pixel_data[38][43] = 0;
        pixel_data[38][44] = 0;
        pixel_data[38][45] = 0;
        pixel_data[38][46] = 0;
        pixel_data[38][47] = 0;
        pixel_data[38][48] = 0;
        pixel_data[38][49] = 0;
        pixel_data[38][50] = 0;
        pixel_data[38][51] = 0;
        pixel_data[38][52] = 0;
        pixel_data[38][53] = 0;
        pixel_data[38][54] = 0;
        pixel_data[38][55] = 0;
        pixel_data[38][56] = 0;
        pixel_data[38][57] = 0;
        pixel_data[38][58] = 0;
        pixel_data[38][59] = 0;
        pixel_data[38][60] = 0;
        pixel_data[38][61] = 0;
        pixel_data[38][62] = 0;
        pixel_data[38][63] = 0;
        pixel_data[38][64] = 0;
        pixel_data[38][65] = 0;
        pixel_data[38][66] = 0;
        pixel_data[38][67] = 0;
        pixel_data[38][68] = 0;
        pixel_data[38][69] = 0;
        pixel_data[38][70] = 0;
        pixel_data[38][71] = 0;
        pixel_data[38][72] = 0;
        pixel_data[38][73] = 0;
        pixel_data[38][74] = 0;
        pixel_data[38][75] = 0;
        pixel_data[38][76] = 0;
        pixel_data[38][77] = 0;
        pixel_data[38][78] = 0;
        pixel_data[38][79] = 0;
        pixel_data[38][80] = 0;
        pixel_data[38][81] = 0;
        pixel_data[38][82] = 0;
        pixel_data[38][83] = 0;
        pixel_data[38][84] = 0;
        pixel_data[38][85] = 0;
        pixel_data[38][86] = 0;
        pixel_data[38][87] = 0;
        pixel_data[38][88] = 0;
        pixel_data[38][89] = 0;
        pixel_data[38][90] = 0;
        pixel_data[38][91] = 0;
        pixel_data[38][92] = 0;
        pixel_data[38][93] = 0;
        pixel_data[38][94] = 0;
        pixel_data[38][95] = 0;
        pixel_data[38][96] = 0;
        pixel_data[38][97] = 0;
        pixel_data[38][98] = 0;
        pixel_data[38][99] = 0;
        pixel_data[38][100] = 0;
        pixel_data[38][101] = 0;
        pixel_data[38][102] = 0;
        pixel_data[38][103] = 0;
        pixel_data[38][104] = 0;
        pixel_data[38][105] = 0;
        pixel_data[38][106] = 0;
        pixel_data[38][107] = 0;
        pixel_data[38][108] = 0;
        pixel_data[38][109] = 0;
        pixel_data[38][110] = 0;
        pixel_data[38][111] = 0;
        pixel_data[38][112] = 0;
        pixel_data[38][113] = 0;
        pixel_data[38][114] = 0;
        pixel_data[38][115] = 0;
        pixel_data[38][116] = 0;
        pixel_data[38][117] = 0;
        pixel_data[38][118] = 0;
        pixel_data[38][119] = 0;
        pixel_data[38][120] = 0;
        pixel_data[38][121] = 0;
        pixel_data[38][122] = 0;
        pixel_data[38][123] = 0;
        pixel_data[38][124] = 0;
        pixel_data[38][125] = 0;
        pixel_data[38][126] = 0;
        pixel_data[38][127] = 0;
        pixel_data[38][128] = 0;
        pixel_data[38][129] = 0;
        pixel_data[38][130] = 0;
        pixel_data[38][131] = 0;
        pixel_data[38][132] = 0;
        pixel_data[38][133] = 0;
        pixel_data[38][134] = 0;
        pixel_data[38][135] = 0;
        pixel_data[38][136] = 0;
        pixel_data[38][137] = 0;
        pixel_data[38][138] = 0;
        pixel_data[38][139] = 0;
        pixel_data[38][140] = 0;
        pixel_data[38][141] = 0;
        pixel_data[38][142] = 0;
        pixel_data[38][143] = 0;
        pixel_data[38][144] = 0;
        pixel_data[38][145] = 0;
        pixel_data[38][146] = 0;
        pixel_data[38][147] = 0;
        pixel_data[38][148] = 0;
        pixel_data[38][149] = 0;
        pixel_data[38][150] = 0;
        pixel_data[38][151] = 0;
        pixel_data[38][152] = 0;
        pixel_data[38][153] = 0;
        pixel_data[38][154] = 0;
        pixel_data[38][155] = 0;
        pixel_data[38][156] = 0;
        pixel_data[38][157] = 0;
        pixel_data[38][158] = 0;
        pixel_data[38][159] = 0;
        pixel_data[38][160] = 0;
        pixel_data[38][161] = 0;
        pixel_data[38][162] = 0;
        pixel_data[38][163] = 0;
        pixel_data[38][164] = 0;
        pixel_data[38][165] = 0;
        pixel_data[38][166] = 0;
        pixel_data[38][167] = 0;
        pixel_data[38][168] = 0;
        pixel_data[38][169] = 0;
        pixel_data[38][170] = 0;
        pixel_data[38][171] = 0;
        pixel_data[38][172] = 0;
        pixel_data[38][173] = 0;
        pixel_data[38][174] = 0;
        pixel_data[38][175] = 0;
        pixel_data[38][176] = 0;
        pixel_data[38][177] = 0;
        pixel_data[38][178] = 0;
        pixel_data[38][179] = 0;
        pixel_data[38][180] = 0;
        pixel_data[38][181] = 0;
        pixel_data[38][182] = 0;
        pixel_data[38][183] = 0;
        pixel_data[38][184] = 0;
        pixel_data[38][185] = 0;
        pixel_data[38][186] = 0;
        pixel_data[38][187] = 0;
        pixel_data[38][188] = 0;
        pixel_data[38][189] = 0;
        pixel_data[38][190] = 0;
        pixel_data[38][191] = 0;
        pixel_data[38][192] = 0;
        pixel_data[38][193] = 0;
        pixel_data[38][194] = 0;
        pixel_data[38][195] = 0;
        pixel_data[38][196] = 0;
        pixel_data[38][197] = 0;
        pixel_data[38][198] = 0;
        pixel_data[38][199] = 0; // y=38
        pixel_data[39][0] = 0;
        pixel_data[39][1] = 0;
        pixel_data[39][2] = 0;
        pixel_data[39][3] = 0;
        pixel_data[39][4] = 0;
        pixel_data[39][5] = 0;
        pixel_data[39][6] = 0;
        pixel_data[39][7] = 0;
        pixel_data[39][8] = 0;
        pixel_data[39][9] = 0;
        pixel_data[39][10] = 0;
        pixel_data[39][11] = 0;
        pixel_data[39][12] = 0;
        pixel_data[39][13] = 0;
        pixel_data[39][14] = 0;
        pixel_data[39][15] = 0;
        pixel_data[39][16] = 0;
        pixel_data[39][17] = 0;
        pixel_data[39][18] = 0;
        pixel_data[39][19] = 0;
        pixel_data[39][20] = 0;
        pixel_data[39][21] = 0;
        pixel_data[39][22] = 0;
        pixel_data[39][23] = 0;
        pixel_data[39][24] = 0;
        pixel_data[39][25] = 0;
        pixel_data[39][26] = 0;
        pixel_data[39][27] = 0;
        pixel_data[39][28] = 0;
        pixel_data[39][29] = 0;
        pixel_data[39][30] = 0;
        pixel_data[39][31] = 0;
        pixel_data[39][32] = 0;
        pixel_data[39][33] = 0;
        pixel_data[39][34] = 0;
        pixel_data[39][35] = 0;
        pixel_data[39][36] = 0;
        pixel_data[39][37] = 0;
        pixel_data[39][38] = 0;
        pixel_data[39][39] = 0;
        pixel_data[39][40] = 0;
        pixel_data[39][41] = 0;
        pixel_data[39][42] = 0;
        pixel_data[39][43] = 0;
        pixel_data[39][44] = 0;
        pixel_data[39][45] = 0;
        pixel_data[39][46] = 0;
        pixel_data[39][47] = 0;
        pixel_data[39][48] = 0;
        pixel_data[39][49] = 0;
        pixel_data[39][50] = 0;
        pixel_data[39][51] = 0;
        pixel_data[39][52] = 0;
        pixel_data[39][53] = 0;
        pixel_data[39][54] = 0;
        pixel_data[39][55] = 0;
        pixel_data[39][56] = 0;
        pixel_data[39][57] = 0;
        pixel_data[39][58] = 0;
        pixel_data[39][59] = 0;
        pixel_data[39][60] = 0;
        pixel_data[39][61] = 0;
        pixel_data[39][62] = 0;
        pixel_data[39][63] = 0;
        pixel_data[39][64] = 0;
        pixel_data[39][65] = 0;
        pixel_data[39][66] = 0;
        pixel_data[39][67] = 0;
        pixel_data[39][68] = 0;
        pixel_data[39][69] = 0;
        pixel_data[39][70] = 0;
        pixel_data[39][71] = 0;
        pixel_data[39][72] = 0;
        pixel_data[39][73] = 0;
        pixel_data[39][74] = 0;
        pixel_data[39][75] = 0;
        pixel_data[39][76] = 0;
        pixel_data[39][77] = 0;
        pixel_data[39][78] = 0;
        pixel_data[39][79] = 0;
        pixel_data[39][80] = 0;
        pixel_data[39][81] = 0;
        pixel_data[39][82] = 0;
        pixel_data[39][83] = 0;
        pixel_data[39][84] = 0;
        pixel_data[39][85] = 0;
        pixel_data[39][86] = 0;
        pixel_data[39][87] = 0;
        pixel_data[39][88] = 0;
        pixel_data[39][89] = 0;
        pixel_data[39][90] = 0;
        pixel_data[39][91] = 0;
        pixel_data[39][92] = 0;
        pixel_data[39][93] = 0;
        pixel_data[39][94] = 0;
        pixel_data[39][95] = 0;
        pixel_data[39][96] = 0;
        pixel_data[39][97] = 0;
        pixel_data[39][98] = 0;
        pixel_data[39][99] = 0;
        pixel_data[39][100] = 0;
        pixel_data[39][101] = 0;
        pixel_data[39][102] = 0;
        pixel_data[39][103] = 0;
        pixel_data[39][104] = 0;
        pixel_data[39][105] = 0;
        pixel_data[39][106] = 0;
        pixel_data[39][107] = 0;
        pixel_data[39][108] = 0;
        pixel_data[39][109] = 0;
        pixel_data[39][110] = 0;
        pixel_data[39][111] = 0;
        pixel_data[39][112] = 0;
        pixel_data[39][113] = 0;
        pixel_data[39][114] = 0;
        pixel_data[39][115] = 0;
        pixel_data[39][116] = 0;
        pixel_data[39][117] = 0;
        pixel_data[39][118] = 0;
        pixel_data[39][119] = 0;
        pixel_data[39][120] = 0;
        pixel_data[39][121] = 0;
        pixel_data[39][122] = 0;
        pixel_data[39][123] = 0;
        pixel_data[39][124] = 0;
        pixel_data[39][125] = 0;
        pixel_data[39][126] = 0;
        pixel_data[39][127] = 0;
        pixel_data[39][128] = 0;
        pixel_data[39][129] = 0;
        pixel_data[39][130] = 0;
        pixel_data[39][131] = 0;
        pixel_data[39][132] = 0;
        pixel_data[39][133] = 0;
        pixel_data[39][134] = 0;
        pixel_data[39][135] = 0;
        pixel_data[39][136] = 0;
        pixel_data[39][137] = 0;
        pixel_data[39][138] = 0;
        pixel_data[39][139] = 0;
        pixel_data[39][140] = 0;
        pixel_data[39][141] = 0;
        pixel_data[39][142] = 0;
        pixel_data[39][143] = 0;
        pixel_data[39][144] = 0;
        pixel_data[39][145] = 0;
        pixel_data[39][146] = 0;
        pixel_data[39][147] = 0;
        pixel_data[39][148] = 0;
        pixel_data[39][149] = 0;
        pixel_data[39][150] = 0;
        pixel_data[39][151] = 0;
        pixel_data[39][152] = 0;
        pixel_data[39][153] = 0;
        pixel_data[39][154] = 0;
        pixel_data[39][155] = 0;
        pixel_data[39][156] = 0;
        pixel_data[39][157] = 0;
        pixel_data[39][158] = 0;
        pixel_data[39][159] = 0;
        pixel_data[39][160] = 0;
        pixel_data[39][161] = 0;
        pixel_data[39][162] = 0;
        pixel_data[39][163] = 0;
        pixel_data[39][164] = 0;
        pixel_data[39][165] = 0;
        pixel_data[39][166] = 0;
        pixel_data[39][167] = 0;
        pixel_data[39][168] = 0;
        pixel_data[39][169] = 0;
        pixel_data[39][170] = 0;
        pixel_data[39][171] = 0;
        pixel_data[39][172] = 0;
        pixel_data[39][173] = 0;
        pixel_data[39][174] = 0;
        pixel_data[39][175] = 0;
        pixel_data[39][176] = 0;
        pixel_data[39][177] = 0;
        pixel_data[39][178] = 0;
        pixel_data[39][179] = 0;
        pixel_data[39][180] = 0;
        pixel_data[39][181] = 0;
        pixel_data[39][182] = 0;
        pixel_data[39][183] = 0;
        pixel_data[39][184] = 0;
        pixel_data[39][185] = 0;
        pixel_data[39][186] = 0;
        pixel_data[39][187] = 0;
        pixel_data[39][188] = 0;
        pixel_data[39][189] = 0;
        pixel_data[39][190] = 0;
        pixel_data[39][191] = 0;
        pixel_data[39][192] = 0;
        pixel_data[39][193] = 0;
        pixel_data[39][194] = 0;
        pixel_data[39][195] = 0;
        pixel_data[39][196] = 0;
        pixel_data[39][197] = 0;
        pixel_data[39][198] = 0;
        pixel_data[39][199] = 0; // y=39
        pixel_data[40][0] = 0;
        pixel_data[40][1] = 0;
        pixel_data[40][2] = 0;
        pixel_data[40][3] = 0;
        pixel_data[40][4] = 0;
        pixel_data[40][5] = 0;
        pixel_data[40][6] = 0;
        pixel_data[40][7] = 0;
        pixel_data[40][8] = 0;
        pixel_data[40][9] = 0;
        pixel_data[40][10] = 0;
        pixel_data[40][11] = 0;
        pixel_data[40][12] = 0;
        pixel_data[40][13] = 0;
        pixel_data[40][14] = 0;
        pixel_data[40][15] = 0;
        pixel_data[40][16] = 0;
        pixel_data[40][17] = 0;
        pixel_data[40][18] = 0;
        pixel_data[40][19] = 0;
        pixel_data[40][20] = 0;
        pixel_data[40][21] = 0;
        pixel_data[40][22] = 0;
        pixel_data[40][23] = 0;
        pixel_data[40][24] = 0;
        pixel_data[40][25] = 0;
        pixel_data[40][26] = 0;
        pixel_data[40][27] = 0;
        pixel_data[40][28] = 0;
        pixel_data[40][29] = 0;
        pixel_data[40][30] = 0;
        pixel_data[40][31] = 0;
        pixel_data[40][32] = 0;
        pixel_data[40][33] = 0;
        pixel_data[40][34] = 0;
        pixel_data[40][35] = 0;
        pixel_data[40][36] = 0;
        pixel_data[40][37] = 0;
        pixel_data[40][38] = 0;
        pixel_data[40][39] = 0;
        pixel_data[40][40] = 0;
        pixel_data[40][41] = 0;
        pixel_data[40][42] = 0;
        pixel_data[40][43] = 0;
        pixel_data[40][44] = 0;
        pixel_data[40][45] = 0;
        pixel_data[40][46] = 0;
        pixel_data[40][47] = 0;
        pixel_data[40][48] = 0;
        pixel_data[40][49] = 0;
        pixel_data[40][50] = 0;
        pixel_data[40][51] = 0;
        pixel_data[40][52] = 0;
        pixel_data[40][53] = 0;
        pixel_data[40][54] = 0;
        pixel_data[40][55] = 0;
        pixel_data[40][56] = 0;
        pixel_data[40][57] = 0;
        pixel_data[40][58] = 0;
        pixel_data[40][59] = 0;
        pixel_data[40][60] = 0;
        pixel_data[40][61] = 0;
        pixel_data[40][62] = 0;
        pixel_data[40][63] = 0;
        pixel_data[40][64] = 0;
        pixel_data[40][65] = 0;
        pixel_data[40][66] = 0;
        pixel_data[40][67] = 0;
        pixel_data[40][68] = 0;
        pixel_data[40][69] = 0;
        pixel_data[40][70] = 0;
        pixel_data[40][71] = 0;
        pixel_data[40][72] = 0;
        pixel_data[40][73] = 0;
        pixel_data[40][74] = 0;
        pixel_data[40][75] = 0;
        pixel_data[40][76] = 0;
        pixel_data[40][77] = 0;
        pixel_data[40][78] = 0;
        pixel_data[40][79] = 0;
        pixel_data[40][80] = 0;
        pixel_data[40][81] = 0;
        pixel_data[40][82] = 0;
        pixel_data[40][83] = 0;
        pixel_data[40][84] = 0;
        pixel_data[40][85] = 0;
        pixel_data[40][86] = 0;
        pixel_data[40][87] = 0;
        pixel_data[40][88] = 0;
        pixel_data[40][89] = 0;
        pixel_data[40][90] = 0;
        pixel_data[40][91] = 0;
        pixel_data[40][92] = 0;
        pixel_data[40][93] = 0;
        pixel_data[40][94] = 0;
        pixel_data[40][95] = 0;
        pixel_data[40][96] = 0;
        pixel_data[40][97] = 0;
        pixel_data[40][98] = 0;
        pixel_data[40][99] = 0;
        pixel_data[40][100] = 0;
        pixel_data[40][101] = 0;
        pixel_data[40][102] = 0;
        pixel_data[40][103] = 0;
        pixel_data[40][104] = 0;
        pixel_data[40][105] = 0;
        pixel_data[40][106] = 0;
        pixel_data[40][107] = 0;
        pixel_data[40][108] = 0;
        pixel_data[40][109] = 0;
        pixel_data[40][110] = 0;
        pixel_data[40][111] = 0;
        pixel_data[40][112] = 0;
        pixel_data[40][113] = 0;
        pixel_data[40][114] = 0;
        pixel_data[40][115] = 0;
        pixel_data[40][116] = 0;
        pixel_data[40][117] = 0;
        pixel_data[40][118] = 0;
        pixel_data[40][119] = 0;
        pixel_data[40][120] = 0;
        pixel_data[40][121] = 0;
        pixel_data[40][122] = 0;
        pixel_data[40][123] = 0;
        pixel_data[40][124] = 0;
        pixel_data[40][125] = 0;
        pixel_data[40][126] = 0;
        pixel_data[40][127] = 0;
        pixel_data[40][128] = 0;
        pixel_data[40][129] = 0;
        pixel_data[40][130] = 0;
        pixel_data[40][131] = 0;
        pixel_data[40][132] = 0;
        pixel_data[40][133] = 0;
        pixel_data[40][134] = 0;
        pixel_data[40][135] = 0;
        pixel_data[40][136] = 0;
        pixel_data[40][137] = 0;
        pixel_data[40][138] = 0;
        pixel_data[40][139] = 0;
        pixel_data[40][140] = 0;
        pixel_data[40][141] = 0;
        pixel_data[40][142] = 0;
        pixel_data[40][143] = 0;
        pixel_data[40][144] = 0;
        pixel_data[40][145] = 0;
        pixel_data[40][146] = 0;
        pixel_data[40][147] = 0;
        pixel_data[40][148] = 0;
        pixel_data[40][149] = 0;
        pixel_data[40][150] = 0;
        pixel_data[40][151] = 0;
        pixel_data[40][152] = 0;
        pixel_data[40][153] = 0;
        pixel_data[40][154] = 0;
        pixel_data[40][155] = 0;
        pixel_data[40][156] = 0;
        pixel_data[40][157] = 0;
        pixel_data[40][158] = 0;
        pixel_data[40][159] = 0;
        pixel_data[40][160] = 0;
        pixel_data[40][161] = 0;
        pixel_data[40][162] = 0;
        pixel_data[40][163] = 0;
        pixel_data[40][164] = 0;
        pixel_data[40][165] = 0;
        pixel_data[40][166] = 0;
        pixel_data[40][167] = 0;
        pixel_data[40][168] = 0;
        pixel_data[40][169] = 0;
        pixel_data[40][170] = 0;
        pixel_data[40][171] = 0;
        pixel_data[40][172] = 0;
        pixel_data[40][173] = 0;
        pixel_data[40][174] = 0;
        pixel_data[40][175] = 0;
        pixel_data[40][176] = 0;
        pixel_data[40][177] = 0;
        pixel_data[40][178] = 0;
        pixel_data[40][179] = 0;
        pixel_data[40][180] = 0;
        pixel_data[40][181] = 0;
        pixel_data[40][182] = 0;
        pixel_data[40][183] = 0;
        pixel_data[40][184] = 0;
        pixel_data[40][185] = 0;
        pixel_data[40][186] = 0;
        pixel_data[40][187] = 0;
        pixel_data[40][188] = 0;
        pixel_data[40][189] = 0;
        pixel_data[40][190] = 0;
        pixel_data[40][191] = 0;
        pixel_data[40][192] = 0;
        pixel_data[40][193] = 0;
        pixel_data[40][194] = 0;
        pixel_data[40][195] = 0;
        pixel_data[40][196] = 0;
        pixel_data[40][197] = 0;
        pixel_data[40][198] = 0;
        pixel_data[40][199] = 0; // y=40
        pixel_data[41][0] = 0;
        pixel_data[41][1] = 0;
        pixel_data[41][2] = 0;
        pixel_data[41][3] = 0;
        pixel_data[41][4] = 0;
        pixel_data[41][5] = 0;
        pixel_data[41][6] = 0;
        pixel_data[41][7] = 0;
        pixel_data[41][8] = 0;
        pixel_data[41][9] = 0;
        pixel_data[41][10] = 0;
        pixel_data[41][11] = 0;
        pixel_data[41][12] = 0;
        pixel_data[41][13] = 0;
        pixel_data[41][14] = 0;
        pixel_data[41][15] = 0;
        pixel_data[41][16] = 0;
        pixel_data[41][17] = 0;
        pixel_data[41][18] = 0;
        pixel_data[41][19] = 0;
        pixel_data[41][20] = 0;
        pixel_data[41][21] = 0;
        pixel_data[41][22] = 0;
        pixel_data[41][23] = 0;
        pixel_data[41][24] = 0;
        pixel_data[41][25] = 0;
        pixel_data[41][26] = 0;
        pixel_data[41][27] = 0;
        pixel_data[41][28] = 0;
        pixel_data[41][29] = 0;
        pixel_data[41][30] = 0;
        pixel_data[41][31] = 0;
        pixel_data[41][32] = 0;
        pixel_data[41][33] = 0;
        pixel_data[41][34] = 0;
        pixel_data[41][35] = 0;
        pixel_data[41][36] = 0;
        pixel_data[41][37] = 0;
        pixel_data[41][38] = 0;
        pixel_data[41][39] = 0;
        pixel_data[41][40] = 0;
        pixel_data[41][41] = 0;
        pixel_data[41][42] = 0;
        pixel_data[41][43] = 0;
        pixel_data[41][44] = 0;
        pixel_data[41][45] = 0;
        pixel_data[41][46] = 0;
        pixel_data[41][47] = 0;
        pixel_data[41][48] = 0;
        pixel_data[41][49] = 0;
        pixel_data[41][50] = 0;
        pixel_data[41][51] = 0;
        pixel_data[41][52] = 0;
        pixel_data[41][53] = 0;
        pixel_data[41][54] = 0;
        pixel_data[41][55] = 0;
        pixel_data[41][56] = 0;
        pixel_data[41][57] = 0;
        pixel_data[41][58] = 0;
        pixel_data[41][59] = 0;
        pixel_data[41][60] = 0;
        pixel_data[41][61] = 0;
        pixel_data[41][62] = 0;
        pixel_data[41][63] = 0;
        pixel_data[41][64] = 0;
        pixel_data[41][65] = 0;
        pixel_data[41][66] = 0;
        pixel_data[41][67] = 0;
        pixel_data[41][68] = 0;
        pixel_data[41][69] = 0;
        pixel_data[41][70] = 0;
        pixel_data[41][71] = 0;
        pixel_data[41][72] = 0;
        pixel_data[41][73] = 0;
        pixel_data[41][74] = 0;
        pixel_data[41][75] = 0;
        pixel_data[41][76] = 0;
        pixel_data[41][77] = 0;
        pixel_data[41][78] = 0;
        pixel_data[41][79] = 0;
        pixel_data[41][80] = 0;
        pixel_data[41][81] = 0;
        pixel_data[41][82] = 0;
        pixel_data[41][83] = 0;
        pixel_data[41][84] = 0;
        pixel_data[41][85] = 0;
        pixel_data[41][86] = 0;
        pixel_data[41][87] = 0;
        pixel_data[41][88] = 0;
        pixel_data[41][89] = 0;
        pixel_data[41][90] = 0;
        pixel_data[41][91] = 0;
        pixel_data[41][92] = 0;
        pixel_data[41][93] = 0;
        pixel_data[41][94] = 0;
        pixel_data[41][95] = 0;
        pixel_data[41][96] = 0;
        pixel_data[41][97] = 0;
        pixel_data[41][98] = 0;
        pixel_data[41][99] = 0;
        pixel_data[41][100] = 0;
        pixel_data[41][101] = 0;
        pixel_data[41][102] = 0;
        pixel_data[41][103] = 0;
        pixel_data[41][104] = 0;
        pixel_data[41][105] = 0;
        pixel_data[41][106] = 0;
        pixel_data[41][107] = 0;
        pixel_data[41][108] = 0;
        pixel_data[41][109] = 0;
        pixel_data[41][110] = 0;
        pixel_data[41][111] = 0;
        pixel_data[41][112] = 0;
        pixel_data[41][113] = 0;
        pixel_data[41][114] = 0;
        pixel_data[41][115] = 0;
        pixel_data[41][116] = 0;
        pixel_data[41][117] = 0;
        pixel_data[41][118] = 0;
        pixel_data[41][119] = 0;
        pixel_data[41][120] = 0;
        pixel_data[41][121] = 0;
        pixel_data[41][122] = 0;
        pixel_data[41][123] = 0;
        pixel_data[41][124] = 0;
        pixel_data[41][125] = 0;
        pixel_data[41][126] = 0;
        pixel_data[41][127] = 0;
        pixel_data[41][128] = 0;
        pixel_data[41][129] = 0;
        pixel_data[41][130] = 0;
        pixel_data[41][131] = 0;
        pixel_data[41][132] = 0;
        pixel_data[41][133] = 0;
        pixel_data[41][134] = 0;
        pixel_data[41][135] = 0;
        pixel_data[41][136] = 0;
        pixel_data[41][137] = 0;
        pixel_data[41][138] = 0;
        pixel_data[41][139] = 0;
        pixel_data[41][140] = 0;
        pixel_data[41][141] = 0;
        pixel_data[41][142] = 0;
        pixel_data[41][143] = 0;
        pixel_data[41][144] = 0;
        pixel_data[41][145] = 0;
        pixel_data[41][146] = 0;
        pixel_data[41][147] = 0;
        pixel_data[41][148] = 0;
        pixel_data[41][149] = 0;
        pixel_data[41][150] = 0;
        pixel_data[41][151] = 0;
        pixel_data[41][152] = 0;
        pixel_data[41][153] = 0;
        pixel_data[41][154] = 0;
        pixel_data[41][155] = 0;
        pixel_data[41][156] = 0;
        pixel_data[41][157] = 0;
        pixel_data[41][158] = 0;
        pixel_data[41][159] = 0;
        pixel_data[41][160] = 0;
        pixel_data[41][161] = 0;
        pixel_data[41][162] = 0;
        pixel_data[41][163] = 0;
        pixel_data[41][164] = 0;
        pixel_data[41][165] = 0;
        pixel_data[41][166] = 0;
        pixel_data[41][167] = 0;
        pixel_data[41][168] = 0;
        pixel_data[41][169] = 0;
        pixel_data[41][170] = 0;
        pixel_data[41][171] = 0;
        pixel_data[41][172] = 0;
        pixel_data[41][173] = 0;
        pixel_data[41][174] = 0;
        pixel_data[41][175] = 0;
        pixel_data[41][176] = 0;
        pixel_data[41][177] = 0;
        pixel_data[41][178] = 0;
        pixel_data[41][179] = 0;
        pixel_data[41][180] = 0;
        pixel_data[41][181] = 0;
        pixel_data[41][182] = 0;
        pixel_data[41][183] = 0;
        pixel_data[41][184] = 0;
        pixel_data[41][185] = 0;
        pixel_data[41][186] = 0;
        pixel_data[41][187] = 0;
        pixel_data[41][188] = 0;
        pixel_data[41][189] = 0;
        pixel_data[41][190] = 0;
        pixel_data[41][191] = 0;
        pixel_data[41][192] = 0;
        pixel_data[41][193] = 0;
        pixel_data[41][194] = 0;
        pixel_data[41][195] = 0;
        pixel_data[41][196] = 0;
        pixel_data[41][197] = 0;
        pixel_data[41][198] = 0;
        pixel_data[41][199] = 0; // y=41
        pixel_data[42][0] = 0;
        pixel_data[42][1] = 0;
        pixel_data[42][2] = 0;
        pixel_data[42][3] = 0;
        pixel_data[42][4] = 0;
        pixel_data[42][5] = 0;
        pixel_data[42][6] = 0;
        pixel_data[42][7] = 0;
        pixel_data[42][8] = 0;
        pixel_data[42][9] = 0;
        pixel_data[42][10] = 0;
        pixel_data[42][11] = 0;
        pixel_data[42][12] = 0;
        pixel_data[42][13] = 0;
        pixel_data[42][14] = 0;
        pixel_data[42][15] = 0;
        pixel_data[42][16] = 0;
        pixel_data[42][17] = 0;
        pixel_data[42][18] = 0;
        pixel_data[42][19] = 0;
        pixel_data[42][20] = 0;
        pixel_data[42][21] = 0;
        pixel_data[42][22] = 0;
        pixel_data[42][23] = 0;
        pixel_data[42][24] = 0;
        pixel_data[42][25] = 0;
        pixel_data[42][26] = 0;
        pixel_data[42][27] = 0;
        pixel_data[42][28] = 0;
        pixel_data[42][29] = 0;
        pixel_data[42][30] = 0;
        pixel_data[42][31] = 0;
        pixel_data[42][32] = 0;
        pixel_data[42][33] = 0;
        pixel_data[42][34] = 0;
        pixel_data[42][35] = 0;
        pixel_data[42][36] = 0;
        pixel_data[42][37] = 0;
        pixel_data[42][38] = 0;
        pixel_data[42][39] = 0;
        pixel_data[42][40] = 0;
        pixel_data[42][41] = 0;
        pixel_data[42][42] = 0;
        pixel_data[42][43] = 0;
        pixel_data[42][44] = 0;
        pixel_data[42][45] = 0;
        pixel_data[42][46] = 0;
        pixel_data[42][47] = 0;
        pixel_data[42][48] = 0;
        pixel_data[42][49] = 0;
        pixel_data[42][50] = 0;
        pixel_data[42][51] = 0;
        pixel_data[42][52] = 0;
        pixel_data[42][53] = 0;
        pixel_data[42][54] = 0;
        pixel_data[42][55] = 0;
        pixel_data[42][56] = 0;
        pixel_data[42][57] = 0;
        pixel_data[42][58] = 0;
        pixel_data[42][59] = 0;
        pixel_data[42][60] = 0;
        pixel_data[42][61] = 0;
        pixel_data[42][62] = 0;
        pixel_data[42][63] = 0;
        pixel_data[42][64] = 0;
        pixel_data[42][65] = 0;
        pixel_data[42][66] = 0;
        pixel_data[42][67] = 0;
        pixel_data[42][68] = 0;
        pixel_data[42][69] = 0;
        pixel_data[42][70] = 0;
        pixel_data[42][71] = 0;
        pixel_data[42][72] = 0;
        pixel_data[42][73] = 0;
        pixel_data[42][74] = 0;
        pixel_data[42][75] = 0;
        pixel_data[42][76] = 0;
        pixel_data[42][77] = 0;
        pixel_data[42][78] = 0;
        pixel_data[42][79] = 0;
        pixel_data[42][80] = 0;
        pixel_data[42][81] = 0;
        pixel_data[42][82] = 0;
        pixel_data[42][83] = 0;
        pixel_data[42][84] = 0;
        pixel_data[42][85] = 0;
        pixel_data[42][86] = 0;
        pixel_data[42][87] = 0;
        pixel_data[42][88] = 0;
        pixel_data[42][89] = 0;
        pixel_data[42][90] = 0;
        pixel_data[42][91] = 0;
        pixel_data[42][92] = 0;
        pixel_data[42][93] = 0;
        pixel_data[42][94] = 0;
        pixel_data[42][95] = 0;
        pixel_data[42][96] = 0;
        pixel_data[42][97] = 0;
        pixel_data[42][98] = 0;
        pixel_data[42][99] = 0;
        pixel_data[42][100] = 0;
        pixel_data[42][101] = 0;
        pixel_data[42][102] = 0;
        pixel_data[42][103] = 0;
        pixel_data[42][104] = 0;
        pixel_data[42][105] = 0;
        pixel_data[42][106] = 0;
        pixel_data[42][107] = 0;
        pixel_data[42][108] = 0;
        pixel_data[42][109] = 0;
        pixel_data[42][110] = 0;
        pixel_data[42][111] = 0;
        pixel_data[42][112] = 0;
        pixel_data[42][113] = 0;
        pixel_data[42][114] = 0;
        pixel_data[42][115] = 0;
        pixel_data[42][116] = 0;
        pixel_data[42][117] = 0;
        pixel_data[42][118] = 0;
        pixel_data[42][119] = 0;
        pixel_data[42][120] = 0;
        pixel_data[42][121] = 0;
        pixel_data[42][122] = 0;
        pixel_data[42][123] = 0;
        pixel_data[42][124] = 0;
        pixel_data[42][125] = 0;
        pixel_data[42][126] = 0;
        pixel_data[42][127] = 0;
        pixel_data[42][128] = 0;
        pixel_data[42][129] = 0;
        pixel_data[42][130] = 0;
        pixel_data[42][131] = 0;
        pixel_data[42][132] = 0;
        pixel_data[42][133] = 0;
        pixel_data[42][134] = 0;
        pixel_data[42][135] = 0;
        pixel_data[42][136] = 0;
        pixel_data[42][137] = 0;
        pixel_data[42][138] = 0;
        pixel_data[42][139] = 0;
        pixel_data[42][140] = 0;
        pixel_data[42][141] = 0;
        pixel_data[42][142] = 0;
        pixel_data[42][143] = 0;
        pixel_data[42][144] = 0;
        pixel_data[42][145] = 0;
        pixel_data[42][146] = 0;
        pixel_data[42][147] = 0;
        pixel_data[42][148] = 0;
        pixel_data[42][149] = 0;
        pixel_data[42][150] = 0;
        pixel_data[42][151] = 0;
        pixel_data[42][152] = 0;
        pixel_data[42][153] = 0;
        pixel_data[42][154] = 0;
        pixel_data[42][155] = 0;
        pixel_data[42][156] = 0;
        pixel_data[42][157] = 0;
        pixel_data[42][158] = 0;
        pixel_data[42][159] = 0;
        pixel_data[42][160] = 0;
        pixel_data[42][161] = 0;
        pixel_data[42][162] = 0;
        pixel_data[42][163] = 0;
        pixel_data[42][164] = 0;
        pixel_data[42][165] = 0;
        pixel_data[42][166] = 0;
        pixel_data[42][167] = 0;
        pixel_data[42][168] = 0;
        pixel_data[42][169] = 0;
        pixel_data[42][170] = 0;
        pixel_data[42][171] = 0;
        pixel_data[42][172] = 0;
        pixel_data[42][173] = 0;
        pixel_data[42][174] = 0;
        pixel_data[42][175] = 0;
        pixel_data[42][176] = 0;
        pixel_data[42][177] = 0;
        pixel_data[42][178] = 0;
        pixel_data[42][179] = 0;
        pixel_data[42][180] = 0;
        pixel_data[42][181] = 0;
        pixel_data[42][182] = 0;
        pixel_data[42][183] = 0;
        pixel_data[42][184] = 0;
        pixel_data[42][185] = 0;
        pixel_data[42][186] = 0;
        pixel_data[42][187] = 0;
        pixel_data[42][188] = 0;
        pixel_data[42][189] = 0;
        pixel_data[42][190] = 0;
        pixel_data[42][191] = 0;
        pixel_data[42][192] = 0;
        pixel_data[42][193] = 0;
        pixel_data[42][194] = 0;
        pixel_data[42][195] = 0;
        pixel_data[42][196] = 0;
        pixel_data[42][197] = 0;
        pixel_data[42][198] = 0;
        pixel_data[42][199] = 0; // y=42
        pixel_data[43][0] = 0;
        pixel_data[43][1] = 0;
        pixel_data[43][2] = 0;
        pixel_data[43][3] = 0;
        pixel_data[43][4] = 0;
        pixel_data[43][5] = 0;
        pixel_data[43][6] = 0;
        pixel_data[43][7] = 0;
        pixel_data[43][8] = 0;
        pixel_data[43][9] = 0;
        pixel_data[43][10] = 0;
        pixel_data[43][11] = 0;
        pixel_data[43][12] = 0;
        pixel_data[43][13] = 0;
        pixel_data[43][14] = 0;
        pixel_data[43][15] = 0;
        pixel_data[43][16] = 0;
        pixel_data[43][17] = 0;
        pixel_data[43][18] = 0;
        pixel_data[43][19] = 0;
        pixel_data[43][20] = 0;
        pixel_data[43][21] = 0;
        pixel_data[43][22] = 0;
        pixel_data[43][23] = 0;
        pixel_data[43][24] = 0;
        pixel_data[43][25] = 0;
        pixel_data[43][26] = 0;
        pixel_data[43][27] = 0;
        pixel_data[43][28] = 0;
        pixel_data[43][29] = 0;
        pixel_data[43][30] = 0;
        pixel_data[43][31] = 0;
        pixel_data[43][32] = 0;
        pixel_data[43][33] = 0;
        pixel_data[43][34] = 0;
        pixel_data[43][35] = 0;
        pixel_data[43][36] = 0;
        pixel_data[43][37] = 0;
        pixel_data[43][38] = 0;
        pixel_data[43][39] = 0;
        pixel_data[43][40] = 0;
        pixel_data[43][41] = 0;
        pixel_data[43][42] = 0;
        pixel_data[43][43] = 0;
        pixel_data[43][44] = 0;
        pixel_data[43][45] = 0;
        pixel_data[43][46] = 0;
        pixel_data[43][47] = 0;
        pixel_data[43][48] = 0;
        pixel_data[43][49] = 0;
        pixel_data[43][50] = 0;
        pixel_data[43][51] = 0;
        pixel_data[43][52] = 0;
        pixel_data[43][53] = 0;
        pixel_data[43][54] = 0;
        pixel_data[43][55] = 0;
        pixel_data[43][56] = 0;
        pixel_data[43][57] = 0;
        pixel_data[43][58] = 0;
        pixel_data[43][59] = 0;
        pixel_data[43][60] = 0;
        pixel_data[43][61] = 0;
        pixel_data[43][62] = 0;
        pixel_data[43][63] = 0;
        pixel_data[43][64] = 0;
        pixel_data[43][65] = 0;
        pixel_data[43][66] = 0;
        pixel_data[43][67] = 0;
        pixel_data[43][68] = 0;
        pixel_data[43][69] = 0;
        pixel_data[43][70] = 0;
        pixel_data[43][71] = 0;
        pixel_data[43][72] = 0;
        pixel_data[43][73] = 0;
        pixel_data[43][74] = 0;
        pixel_data[43][75] = 0;
        pixel_data[43][76] = 0;
        pixel_data[43][77] = 0;
        pixel_data[43][78] = 0;
        pixel_data[43][79] = 0;
        pixel_data[43][80] = 0;
        pixel_data[43][81] = 0;
        pixel_data[43][82] = 0;
        pixel_data[43][83] = 0;
        pixel_data[43][84] = 0;
        pixel_data[43][85] = 0;
        pixel_data[43][86] = 0;
        pixel_data[43][87] = 0;
        pixel_data[43][88] = 0;
        pixel_data[43][89] = 0;
        pixel_data[43][90] = 0;
        pixel_data[43][91] = 0;
        pixel_data[43][92] = 0;
        pixel_data[43][93] = 0;
        pixel_data[43][94] = 0;
        pixel_data[43][95] = 0;
        pixel_data[43][96] = 0;
        pixel_data[43][97] = 0;
        pixel_data[43][98] = 0;
        pixel_data[43][99] = 0;
        pixel_data[43][100] = 0;
        pixel_data[43][101] = 0;
        pixel_data[43][102] = 0;
        pixel_data[43][103] = 0;
        pixel_data[43][104] = 0;
        pixel_data[43][105] = 0;
        pixel_data[43][106] = 0;
        pixel_data[43][107] = 0;
        pixel_data[43][108] = 0;
        pixel_data[43][109] = 0;
        pixel_data[43][110] = 0;
        pixel_data[43][111] = 0;
        pixel_data[43][112] = 0;
        pixel_data[43][113] = 0;
        pixel_data[43][114] = 0;
        pixel_data[43][115] = 0;
        pixel_data[43][116] = 0;
        pixel_data[43][117] = 0;
        pixel_data[43][118] = 0;
        pixel_data[43][119] = 0;
        pixel_data[43][120] = 0;
        pixel_data[43][121] = 0;
        pixel_data[43][122] = 0;
        pixel_data[43][123] = 0;
        pixel_data[43][124] = 0;
        pixel_data[43][125] = 0;
        pixel_data[43][126] = 0;
        pixel_data[43][127] = 0;
        pixel_data[43][128] = 0;
        pixel_data[43][129] = 0;
        pixel_data[43][130] = 0;
        pixel_data[43][131] = 0;
        pixel_data[43][132] = 0;
        pixel_data[43][133] = 0;
        pixel_data[43][134] = 0;
        pixel_data[43][135] = 0;
        pixel_data[43][136] = 0;
        pixel_data[43][137] = 0;
        pixel_data[43][138] = 0;
        pixel_data[43][139] = 0;
        pixel_data[43][140] = 0;
        pixel_data[43][141] = 0;
        pixel_data[43][142] = 0;
        pixel_data[43][143] = 0;
        pixel_data[43][144] = 0;
        pixel_data[43][145] = 0;
        pixel_data[43][146] = 0;
        pixel_data[43][147] = 0;
        pixel_data[43][148] = 0;
        pixel_data[43][149] = 0;
        pixel_data[43][150] = 0;
        pixel_data[43][151] = 0;
        pixel_data[43][152] = 0;
        pixel_data[43][153] = 0;
        pixel_data[43][154] = 0;
        pixel_data[43][155] = 0;
        pixel_data[43][156] = 0;
        pixel_data[43][157] = 0;
        pixel_data[43][158] = 0;
        pixel_data[43][159] = 0;
        pixel_data[43][160] = 0;
        pixel_data[43][161] = 0;
        pixel_data[43][162] = 0;
        pixel_data[43][163] = 0;
        pixel_data[43][164] = 0;
        pixel_data[43][165] = 0;
        pixel_data[43][166] = 0;
        pixel_data[43][167] = 0;
        pixel_data[43][168] = 0;
        pixel_data[43][169] = 0;
        pixel_data[43][170] = 0;
        pixel_data[43][171] = 0;
        pixel_data[43][172] = 0;
        pixel_data[43][173] = 0;
        pixel_data[43][174] = 0;
        pixel_data[43][175] = 0;
        pixel_data[43][176] = 0;
        pixel_data[43][177] = 0;
        pixel_data[43][178] = 0;
        pixel_data[43][179] = 0;
        pixel_data[43][180] = 0;
        pixel_data[43][181] = 0;
        pixel_data[43][182] = 0;
        pixel_data[43][183] = 0;
        pixel_data[43][184] = 0;
        pixel_data[43][185] = 0;
        pixel_data[43][186] = 0;
        pixel_data[43][187] = 0;
        pixel_data[43][188] = 0;
        pixel_data[43][189] = 0;
        pixel_data[43][190] = 0;
        pixel_data[43][191] = 0;
        pixel_data[43][192] = 0;
        pixel_data[43][193] = 0;
        pixel_data[43][194] = 0;
        pixel_data[43][195] = 0;
        pixel_data[43][196] = 0;
        pixel_data[43][197] = 0;
        pixel_data[43][198] = 0;
        pixel_data[43][199] = 0; // y=43
        pixel_data[44][0] = 0;
        pixel_data[44][1] = 0;
        pixel_data[44][2] = 0;
        pixel_data[44][3] = 0;
        pixel_data[44][4] = 0;
        pixel_data[44][5] = 0;
        pixel_data[44][6] = 0;
        pixel_data[44][7] = 0;
        pixel_data[44][8] = 0;
        pixel_data[44][9] = 0;
        pixel_data[44][10] = 0;
        pixel_data[44][11] = 0;
        pixel_data[44][12] = 0;
        pixel_data[44][13] = 0;
        pixel_data[44][14] = 0;
        pixel_data[44][15] = 0;
        pixel_data[44][16] = 0;
        pixel_data[44][17] = 0;
        pixel_data[44][18] = 0;
        pixel_data[44][19] = 0;
        pixel_data[44][20] = 0;
        pixel_data[44][21] = 0;
        pixel_data[44][22] = 0;
        pixel_data[44][23] = 0;
        pixel_data[44][24] = 0;
        pixel_data[44][25] = 0;
        pixel_data[44][26] = 0;
        pixel_data[44][27] = 0;
        pixel_data[44][28] = 0;
        pixel_data[44][29] = 0;
        pixel_data[44][30] = 0;
        pixel_data[44][31] = 0;
        pixel_data[44][32] = 0;
        pixel_data[44][33] = 0;
        pixel_data[44][34] = 0;
        pixel_data[44][35] = 0;
        pixel_data[44][36] = 0;
        pixel_data[44][37] = 0;
        pixel_data[44][38] = 0;
        pixel_data[44][39] = 0;
        pixel_data[44][40] = 0;
        pixel_data[44][41] = 0;
        pixel_data[44][42] = 0;
        pixel_data[44][43] = 0;
        pixel_data[44][44] = 0;
        pixel_data[44][45] = 0;
        pixel_data[44][46] = 0;
        pixel_data[44][47] = 0;
        pixel_data[44][48] = 0;
        pixel_data[44][49] = 0;
        pixel_data[44][50] = 0;
        pixel_data[44][51] = 0;
        pixel_data[44][52] = 0;
        pixel_data[44][53] = 0;
        pixel_data[44][54] = 0;
        pixel_data[44][55] = 0;
        pixel_data[44][56] = 0;
        pixel_data[44][57] = 0;
        pixel_data[44][58] = 0;
        pixel_data[44][59] = 0;
        pixel_data[44][60] = 0;
        pixel_data[44][61] = 0;
        pixel_data[44][62] = 0;
        pixel_data[44][63] = 0;
        pixel_data[44][64] = 0;
        pixel_data[44][65] = 0;
        pixel_data[44][66] = 0;
        pixel_data[44][67] = 0;
        pixel_data[44][68] = 0;
        pixel_data[44][69] = 0;
        pixel_data[44][70] = 0;
        pixel_data[44][71] = 0;
        pixel_data[44][72] = 0;
        pixel_data[44][73] = 0;
        pixel_data[44][74] = 0;
        pixel_data[44][75] = 0;
        pixel_data[44][76] = 0;
        pixel_data[44][77] = 0;
        pixel_data[44][78] = 0;
        pixel_data[44][79] = 0;
        pixel_data[44][80] = 0;
        pixel_data[44][81] = 0;
        pixel_data[44][82] = 0;
        pixel_data[44][83] = 0;
        pixel_data[44][84] = 0;
        pixel_data[44][85] = 0;
        pixel_data[44][86] = 0;
        pixel_data[44][87] = 0;
        pixel_data[44][88] = 0;
        pixel_data[44][89] = 0;
        pixel_data[44][90] = 0;
        pixel_data[44][91] = 0;
        pixel_data[44][92] = 0;
        pixel_data[44][93] = 0;
        pixel_data[44][94] = 0;
        pixel_data[44][95] = 0;
        pixel_data[44][96] = 0;
        pixel_data[44][97] = 0;
        pixel_data[44][98] = 0;
        pixel_data[44][99] = 0;
        pixel_data[44][100] = 0;
        pixel_data[44][101] = 0;
        pixel_data[44][102] = 0;
        pixel_data[44][103] = 0;
        pixel_data[44][104] = 0;
        pixel_data[44][105] = 0;
        pixel_data[44][106] = 0;
        pixel_data[44][107] = 0;
        pixel_data[44][108] = 0;
        pixel_data[44][109] = 0;
        pixel_data[44][110] = 0;
        pixel_data[44][111] = 0;
        pixel_data[44][112] = 0;
        pixel_data[44][113] = 0;
        pixel_data[44][114] = 0;
        pixel_data[44][115] = 0;
        pixel_data[44][116] = 0;
        pixel_data[44][117] = 0;
        pixel_data[44][118] = 0;
        pixel_data[44][119] = 0;
        pixel_data[44][120] = 0;
        pixel_data[44][121] = 0;
        pixel_data[44][122] = 0;
        pixel_data[44][123] = 0;
        pixel_data[44][124] = 0;
        pixel_data[44][125] = 0;
        pixel_data[44][126] = 0;
        pixel_data[44][127] = 0;
        pixel_data[44][128] = 0;
        pixel_data[44][129] = 0;
        pixel_data[44][130] = 0;
        pixel_data[44][131] = 0;
        pixel_data[44][132] = 0;
        pixel_data[44][133] = 0;
        pixel_data[44][134] = 0;
        pixel_data[44][135] = 0;
        pixel_data[44][136] = 0;
        pixel_data[44][137] = 0;
        pixel_data[44][138] = 0;
        pixel_data[44][139] = 0;
        pixel_data[44][140] = 0;
        pixel_data[44][141] = 0;
        pixel_data[44][142] = 0;
        pixel_data[44][143] = 0;
        pixel_data[44][144] = 0;
        pixel_data[44][145] = 0;
        pixel_data[44][146] = 0;
        pixel_data[44][147] = 0;
        pixel_data[44][148] = 0;
        pixel_data[44][149] = 0;
        pixel_data[44][150] = 0;
        pixel_data[44][151] = 0;
        pixel_data[44][152] = 0;
        pixel_data[44][153] = 0;
        pixel_data[44][154] = 0;
        pixel_data[44][155] = 0;
        pixel_data[44][156] = 0;
        pixel_data[44][157] = 0;
        pixel_data[44][158] = 0;
        pixel_data[44][159] = 0;
        pixel_data[44][160] = 0;
        pixel_data[44][161] = 0;
        pixel_data[44][162] = 0;
        pixel_data[44][163] = 0;
        pixel_data[44][164] = 0;
        pixel_data[44][165] = 0;
        pixel_data[44][166] = 0;
        pixel_data[44][167] = 0;
        pixel_data[44][168] = 0;
        pixel_data[44][169] = 0;
        pixel_data[44][170] = 0;
        pixel_data[44][171] = 0;
        pixel_data[44][172] = 0;
        pixel_data[44][173] = 0;
        pixel_data[44][174] = 0;
        pixel_data[44][175] = 0;
        pixel_data[44][176] = 0;
        pixel_data[44][177] = 0;
        pixel_data[44][178] = 0;
        pixel_data[44][179] = 0;
        pixel_data[44][180] = 0;
        pixel_data[44][181] = 0;
        pixel_data[44][182] = 0;
        pixel_data[44][183] = 0;
        pixel_data[44][184] = 0;
        pixel_data[44][185] = 0;
        pixel_data[44][186] = 0;
        pixel_data[44][187] = 0;
        pixel_data[44][188] = 0;
        pixel_data[44][189] = 0;
        pixel_data[44][190] = 0;
        pixel_data[44][191] = 0;
        pixel_data[44][192] = 0;
        pixel_data[44][193] = 0;
        pixel_data[44][194] = 0;
        pixel_data[44][195] = 0;
        pixel_data[44][196] = 0;
        pixel_data[44][197] = 0;
        pixel_data[44][198] = 0;
        pixel_data[44][199] = 0; // y=44
        pixel_data[45][0] = 0;
        pixel_data[45][1] = 0;
        pixel_data[45][2] = 0;
        pixel_data[45][3] = 0;
        pixel_data[45][4] = 0;
        pixel_data[45][5] = 0;
        pixel_data[45][6] = 0;
        pixel_data[45][7] = 0;
        pixel_data[45][8] = 0;
        pixel_data[45][9] = 0;
        pixel_data[45][10] = 0;
        pixel_data[45][11] = 0;
        pixel_data[45][12] = 0;
        pixel_data[45][13] = 0;
        pixel_data[45][14] = 0;
        pixel_data[45][15] = 0;
        pixel_data[45][16] = 0;
        pixel_data[45][17] = 0;
        pixel_data[45][18] = 0;
        pixel_data[45][19] = 0;
        pixel_data[45][20] = 0;
        pixel_data[45][21] = 0;
        pixel_data[45][22] = 0;
        pixel_data[45][23] = 0;
        pixel_data[45][24] = 0;
        pixel_data[45][25] = 0;
        pixel_data[45][26] = 0;
        pixel_data[45][27] = 0;
        pixel_data[45][28] = 0;
        pixel_data[45][29] = 0;
        pixel_data[45][30] = 0;
        pixel_data[45][31] = 0;
        pixel_data[45][32] = 0;
        pixel_data[45][33] = 0;
        pixel_data[45][34] = 0;
        pixel_data[45][35] = 0;
        pixel_data[45][36] = 0;
        pixel_data[45][37] = 0;
        pixel_data[45][38] = 0;
        pixel_data[45][39] = 0;
        pixel_data[45][40] = 0;
        pixel_data[45][41] = 0;
        pixel_data[45][42] = 0;
        pixel_data[45][43] = 0;
        pixel_data[45][44] = 0;
        pixel_data[45][45] = 0;
        pixel_data[45][46] = 0;
        pixel_data[45][47] = 0;
        pixel_data[45][48] = 0;
        pixel_data[45][49] = 0;
        pixel_data[45][50] = 0;
        pixel_data[45][51] = 0;
        pixel_data[45][52] = 0;
        pixel_data[45][53] = 0;
        pixel_data[45][54] = 0;
        pixel_data[45][55] = 0;
        pixel_data[45][56] = 0;
        pixel_data[45][57] = 0;
        pixel_data[45][58] = 0;
        pixel_data[45][59] = 0;
        pixel_data[45][60] = 0;
        pixel_data[45][61] = 0;
        pixel_data[45][62] = 0;
        pixel_data[45][63] = 0;
        pixel_data[45][64] = 0;
        pixel_data[45][65] = 0;
        pixel_data[45][66] = 0;
        pixel_data[45][67] = 0;
        pixel_data[45][68] = 0;
        pixel_data[45][69] = 0;
        pixel_data[45][70] = 0;
        pixel_data[45][71] = 0;
        pixel_data[45][72] = 0;
        pixel_data[45][73] = 0;
        pixel_data[45][74] = 0;
        pixel_data[45][75] = 0;
        pixel_data[45][76] = 0;
        pixel_data[45][77] = 0;
        pixel_data[45][78] = 0;
        pixel_data[45][79] = 0;
        pixel_data[45][80] = 0;
        pixel_data[45][81] = 0;
        pixel_data[45][82] = 0;
        pixel_data[45][83] = 0;
        pixel_data[45][84] = 0;
        pixel_data[45][85] = 0;
        pixel_data[45][86] = 0;
        pixel_data[45][87] = 0;
        pixel_data[45][88] = 0;
        pixel_data[45][89] = 0;
        pixel_data[45][90] = 0;
        pixel_data[45][91] = 0;
        pixel_data[45][92] = 0;
        pixel_data[45][93] = 0;
        pixel_data[45][94] = 0;
        pixel_data[45][95] = 0;
        pixel_data[45][96] = 0;
        pixel_data[45][97] = 0;
        pixel_data[45][98] = 0;
        pixel_data[45][99] = 0;
        pixel_data[45][100] = 0;
        pixel_data[45][101] = 0;
        pixel_data[45][102] = 0;
        pixel_data[45][103] = 0;
        pixel_data[45][104] = 0;
        pixel_data[45][105] = 0;
        pixel_data[45][106] = 0;
        pixel_data[45][107] = 0;
        pixel_data[45][108] = 0;
        pixel_data[45][109] = 0;
        pixel_data[45][110] = 0;
        pixel_data[45][111] = 0;
        pixel_data[45][112] = 0;
        pixel_data[45][113] = 0;
        pixel_data[45][114] = 0;
        pixel_data[45][115] = 0;
        pixel_data[45][116] = 0;
        pixel_data[45][117] = 0;
        pixel_data[45][118] = 0;
        pixel_data[45][119] = 0;
        pixel_data[45][120] = 0;
        pixel_data[45][121] = 0;
        pixel_data[45][122] = 0;
        pixel_data[45][123] = 0;
        pixel_data[45][124] = 0;
        pixel_data[45][125] = 0;
        pixel_data[45][126] = 0;
        pixel_data[45][127] = 0;
        pixel_data[45][128] = 0;
        pixel_data[45][129] = 0;
        pixel_data[45][130] = 0;
        pixel_data[45][131] = 0;
        pixel_data[45][132] = 0;
        pixel_data[45][133] = 0;
        pixel_data[45][134] = 0;
        pixel_data[45][135] = 0;
        pixel_data[45][136] = 0;
        pixel_data[45][137] = 0;
        pixel_data[45][138] = 0;
        pixel_data[45][139] = 0;
        pixel_data[45][140] = 0;
        pixel_data[45][141] = 0;
        pixel_data[45][142] = 0;
        pixel_data[45][143] = 0;
        pixel_data[45][144] = 0;
        pixel_data[45][145] = 0;
        pixel_data[45][146] = 0;
        pixel_data[45][147] = 0;
        pixel_data[45][148] = 0;
        pixel_data[45][149] = 0;
        pixel_data[45][150] = 0;
        pixel_data[45][151] = 0;
        pixel_data[45][152] = 0;
        pixel_data[45][153] = 0;
        pixel_data[45][154] = 0;
        pixel_data[45][155] = 0;
        pixel_data[45][156] = 0;
        pixel_data[45][157] = 0;
        pixel_data[45][158] = 0;
        pixel_data[45][159] = 0;
        pixel_data[45][160] = 0;
        pixel_data[45][161] = 0;
        pixel_data[45][162] = 0;
        pixel_data[45][163] = 0;
        pixel_data[45][164] = 0;
        pixel_data[45][165] = 0;
        pixel_data[45][166] = 0;
        pixel_data[45][167] = 0;
        pixel_data[45][168] = 0;
        pixel_data[45][169] = 0;
        pixel_data[45][170] = 0;
        pixel_data[45][171] = 0;
        pixel_data[45][172] = 0;
        pixel_data[45][173] = 0;
        pixel_data[45][174] = 0;
        pixel_data[45][175] = 0;
        pixel_data[45][176] = 0;
        pixel_data[45][177] = 0;
        pixel_data[45][178] = 0;
        pixel_data[45][179] = 0;
        pixel_data[45][180] = 0;
        pixel_data[45][181] = 0;
        pixel_data[45][182] = 0;
        pixel_data[45][183] = 0;
        pixel_data[45][184] = 0;
        pixel_data[45][185] = 0;
        pixel_data[45][186] = 0;
        pixel_data[45][187] = 0;
        pixel_data[45][188] = 0;
        pixel_data[45][189] = 0;
        pixel_data[45][190] = 0;
        pixel_data[45][191] = 0;
        pixel_data[45][192] = 0;
        pixel_data[45][193] = 0;
        pixel_data[45][194] = 0;
        pixel_data[45][195] = 0;
        pixel_data[45][196] = 0;
        pixel_data[45][197] = 0;
        pixel_data[45][198] = 0;
        pixel_data[45][199] = 0; // y=45
        pixel_data[46][0] = 0;
        pixel_data[46][1] = 0;
        pixel_data[46][2] = 0;
        pixel_data[46][3] = 0;
        pixel_data[46][4] = 0;
        pixel_data[46][5] = 0;
        pixel_data[46][6] = 0;
        pixel_data[46][7] = 0;
        pixel_data[46][8] = 0;
        pixel_data[46][9] = 0;
        pixel_data[46][10] = 0;
        pixel_data[46][11] = 0;
        pixel_data[46][12] = 0;
        pixel_data[46][13] = 0;
        pixel_data[46][14] = 0;
        pixel_data[46][15] = 0;
        pixel_data[46][16] = 0;
        pixel_data[46][17] = 0;
        pixel_data[46][18] = 0;
        pixel_data[46][19] = 0;
        pixel_data[46][20] = 0;
        pixel_data[46][21] = 0;
        pixel_data[46][22] = 0;
        pixel_data[46][23] = 0;
        pixel_data[46][24] = 0;
        pixel_data[46][25] = 0;
        pixel_data[46][26] = 0;
        pixel_data[46][27] = 0;
        pixel_data[46][28] = 0;
        pixel_data[46][29] = 0;
        pixel_data[46][30] = 0;
        pixel_data[46][31] = 0;
        pixel_data[46][32] = 0;
        pixel_data[46][33] = 0;
        pixel_data[46][34] = 0;
        pixel_data[46][35] = 0;
        pixel_data[46][36] = 0;
        pixel_data[46][37] = 0;
        pixel_data[46][38] = 0;
        pixel_data[46][39] = 0;
        pixel_data[46][40] = 0;
        pixel_data[46][41] = 0;
        pixel_data[46][42] = 0;
        pixel_data[46][43] = 0;
        pixel_data[46][44] = 0;
        pixel_data[46][45] = 0;
        pixel_data[46][46] = 0;
        pixel_data[46][47] = 0;
        pixel_data[46][48] = 0;
        pixel_data[46][49] = 0;
        pixel_data[46][50] = 0;
        pixel_data[46][51] = 0;
        pixel_data[46][52] = 0;
        pixel_data[46][53] = 0;
        pixel_data[46][54] = 0;
        pixel_data[46][55] = 0;
        pixel_data[46][56] = 0;
        pixel_data[46][57] = 0;
        pixel_data[46][58] = 0;
        pixel_data[46][59] = 0;
        pixel_data[46][60] = 0;
        pixel_data[46][61] = 0;
        pixel_data[46][62] = 0;
        pixel_data[46][63] = 0;
        pixel_data[46][64] = 0;
        pixel_data[46][65] = 0;
        pixel_data[46][66] = 0;
        pixel_data[46][67] = 0;
        pixel_data[46][68] = 0;
        pixel_data[46][69] = 0;
        pixel_data[46][70] = 0;
        pixel_data[46][71] = 0;
        pixel_data[46][72] = 0;
        pixel_data[46][73] = 0;
        pixel_data[46][74] = 0;
        pixel_data[46][75] = 0;
        pixel_data[46][76] = 0;
        pixel_data[46][77] = 0;
        pixel_data[46][78] = 0;
        pixel_data[46][79] = 0;
        pixel_data[46][80] = 0;
        pixel_data[46][81] = 0;
        pixel_data[46][82] = 0;
        pixel_data[46][83] = 0;
        pixel_data[46][84] = 0;
        pixel_data[46][85] = 0;
        pixel_data[46][86] = 0;
        pixel_data[46][87] = 0;
        pixel_data[46][88] = 0;
        pixel_data[46][89] = 0;
        pixel_data[46][90] = 0;
        pixel_data[46][91] = 0;
        pixel_data[46][92] = 0;
        pixel_data[46][93] = 0;
        pixel_data[46][94] = 0;
        pixel_data[46][95] = 0;
        pixel_data[46][96] = 0;
        pixel_data[46][97] = 0;
        pixel_data[46][98] = 0;
        pixel_data[46][99] = 0;
        pixel_data[46][100] = 0;
        pixel_data[46][101] = 0;
        pixel_data[46][102] = 0;
        pixel_data[46][103] = 0;
        pixel_data[46][104] = 0;
        pixel_data[46][105] = 0;
        pixel_data[46][106] = 0;
        pixel_data[46][107] = 0;
        pixel_data[46][108] = 0;
        pixel_data[46][109] = 0;
        pixel_data[46][110] = 0;
        pixel_data[46][111] = 0;
        pixel_data[46][112] = 0;
        pixel_data[46][113] = 0;
        pixel_data[46][114] = 0;
        pixel_data[46][115] = 0;
        pixel_data[46][116] = 0;
        pixel_data[46][117] = 0;
        pixel_data[46][118] = 0;
        pixel_data[46][119] = 0;
        pixel_data[46][120] = 0;
        pixel_data[46][121] = 0;
        pixel_data[46][122] = 0;
        pixel_data[46][123] = 0;
        pixel_data[46][124] = 0;
        pixel_data[46][125] = 0;
        pixel_data[46][126] = 0;
        pixel_data[46][127] = 0;
        pixel_data[46][128] = 0;
        pixel_data[46][129] = 0;
        pixel_data[46][130] = 0;
        pixel_data[46][131] = 0;
        pixel_data[46][132] = 0;
        pixel_data[46][133] = 0;
        pixel_data[46][134] = 0;
        pixel_data[46][135] = 0;
        pixel_data[46][136] = 0;
        pixel_data[46][137] = 0;
        pixel_data[46][138] = 0;
        pixel_data[46][139] = 0;
        pixel_data[46][140] = 0;
        pixel_data[46][141] = 0;
        pixel_data[46][142] = 0;
        pixel_data[46][143] = 0;
        pixel_data[46][144] = 0;
        pixel_data[46][145] = 0;
        pixel_data[46][146] = 0;
        pixel_data[46][147] = 0;
        pixel_data[46][148] = 0;
        pixel_data[46][149] = 0;
        pixel_data[46][150] = 0;
        pixel_data[46][151] = 0;
        pixel_data[46][152] = 0;
        pixel_data[46][153] = 0;
        pixel_data[46][154] = 0;
        pixel_data[46][155] = 0;
        pixel_data[46][156] = 0;
        pixel_data[46][157] = 0;
        pixel_data[46][158] = 0;
        pixel_data[46][159] = 0;
        pixel_data[46][160] = 0;
        pixel_data[46][161] = 0;
        pixel_data[46][162] = 0;
        pixel_data[46][163] = 0;
        pixel_data[46][164] = 0;
        pixel_data[46][165] = 0;
        pixel_data[46][166] = 0;
        pixel_data[46][167] = 0;
        pixel_data[46][168] = 0;
        pixel_data[46][169] = 0;
        pixel_data[46][170] = 0;
        pixel_data[46][171] = 0;
        pixel_data[46][172] = 0;
        pixel_data[46][173] = 0;
        pixel_data[46][174] = 0;
        pixel_data[46][175] = 0;
        pixel_data[46][176] = 0;
        pixel_data[46][177] = 0;
        pixel_data[46][178] = 0;
        pixel_data[46][179] = 0;
        pixel_data[46][180] = 0;
        pixel_data[46][181] = 0;
        pixel_data[46][182] = 0;
        pixel_data[46][183] = 0;
        pixel_data[46][184] = 0;
        pixel_data[46][185] = 0;
        pixel_data[46][186] = 0;
        pixel_data[46][187] = 0;
        pixel_data[46][188] = 0;
        pixel_data[46][189] = 0;
        pixel_data[46][190] = 0;
        pixel_data[46][191] = 0;
        pixel_data[46][192] = 0;
        pixel_data[46][193] = 0;
        pixel_data[46][194] = 0;
        pixel_data[46][195] = 0;
        pixel_data[46][196] = 0;
        pixel_data[46][197] = 0;
        pixel_data[46][198] = 0;
        pixel_data[46][199] = 0; // y=46
        pixel_data[47][0] = 0;
        pixel_data[47][1] = 0;
        pixel_data[47][2] = 0;
        pixel_data[47][3] = 0;
        pixel_data[47][4] = 0;
        pixel_data[47][5] = 0;
        pixel_data[47][6] = 0;
        pixel_data[47][7] = 0;
        pixel_data[47][8] = 0;
        pixel_data[47][9] = 0;
        pixel_data[47][10] = 0;
        pixel_data[47][11] = 0;
        pixel_data[47][12] = 0;
        pixel_data[47][13] = 0;
        pixel_data[47][14] = 0;
        pixel_data[47][15] = 0;
        pixel_data[47][16] = 0;
        pixel_data[47][17] = 0;
        pixel_data[47][18] = 0;
        pixel_data[47][19] = 0;
        pixel_data[47][20] = 0;
        pixel_data[47][21] = 0;
        pixel_data[47][22] = 0;
        pixel_data[47][23] = 0;
        pixel_data[47][24] = 0;
        pixel_data[47][25] = 0;
        pixel_data[47][26] = 0;
        pixel_data[47][27] = 0;
        pixel_data[47][28] = 0;
        pixel_data[47][29] = 0;
        pixel_data[47][30] = 0;
        pixel_data[47][31] = 0;
        pixel_data[47][32] = 0;
        pixel_data[47][33] = 0;
        pixel_data[47][34] = 0;
        pixel_data[47][35] = 0;
        pixel_data[47][36] = 0;
        pixel_data[47][37] = 0;
        pixel_data[47][38] = 0;
        pixel_data[47][39] = 0;
        pixel_data[47][40] = 0;
        pixel_data[47][41] = 0;
        pixel_data[47][42] = 0;
        pixel_data[47][43] = 0;
        pixel_data[47][44] = 0;
        pixel_data[47][45] = 0;
        pixel_data[47][46] = 0;
        pixel_data[47][47] = 0;
        pixel_data[47][48] = 0;
        pixel_data[47][49] = 0;
        pixel_data[47][50] = 0;
        pixel_data[47][51] = 0;
        pixel_data[47][52] = 0;
        pixel_data[47][53] = 0;
        pixel_data[47][54] = 0;
        pixel_data[47][55] = 0;
        pixel_data[47][56] = 0;
        pixel_data[47][57] = 0;
        pixel_data[47][58] = 0;
        pixel_data[47][59] = 0;
        pixel_data[47][60] = 0;
        pixel_data[47][61] = 0;
        pixel_data[47][62] = 0;
        pixel_data[47][63] = 0;
        pixel_data[47][64] = 0;
        pixel_data[47][65] = 0;
        pixel_data[47][66] = 0;
        pixel_data[47][67] = 0;
        pixel_data[47][68] = 0;
        pixel_data[47][69] = 0;
        pixel_data[47][70] = 0;
        pixel_data[47][71] = 0;
        pixel_data[47][72] = 0;
        pixel_data[47][73] = 0;
        pixel_data[47][74] = 0;
        pixel_data[47][75] = 0;
        pixel_data[47][76] = 0;
        pixel_data[47][77] = 0;
        pixel_data[47][78] = 0;
        pixel_data[47][79] = 0;
        pixel_data[47][80] = 0;
        pixel_data[47][81] = 0;
        pixel_data[47][82] = 0;
        pixel_data[47][83] = 0;
        pixel_data[47][84] = 0;
        pixel_data[47][85] = 0;
        pixel_data[47][86] = 0;
        pixel_data[47][87] = 0;
        pixel_data[47][88] = 0;
        pixel_data[47][89] = 0;
        pixel_data[47][90] = 0;
        pixel_data[47][91] = 0;
        pixel_data[47][92] = 0;
        pixel_data[47][93] = 0;
        pixel_data[47][94] = 0;
        pixel_data[47][95] = 0;
        pixel_data[47][96] = 0;
        pixel_data[47][97] = 0;
        pixel_data[47][98] = 0;
        pixel_data[47][99] = 0;
        pixel_data[47][100] = 0;
        pixel_data[47][101] = 0;
        pixel_data[47][102] = 0;
        pixel_data[47][103] = 0;
        pixel_data[47][104] = 0;
        pixel_data[47][105] = 0;
        pixel_data[47][106] = 0;
        pixel_data[47][107] = 0;
        pixel_data[47][108] = 0;
        pixel_data[47][109] = 0;
        pixel_data[47][110] = 0;
        pixel_data[47][111] = 0;
        pixel_data[47][112] = 0;
        pixel_data[47][113] = 0;
        pixel_data[47][114] = 0;
        pixel_data[47][115] = 0;
        pixel_data[47][116] = 0;
        pixel_data[47][117] = 0;
        pixel_data[47][118] = 0;
        pixel_data[47][119] = 0;
        pixel_data[47][120] = 0;
        pixel_data[47][121] = 0;
        pixel_data[47][122] = 0;
        pixel_data[47][123] = 0;
        pixel_data[47][124] = 0;
        pixel_data[47][125] = 0;
        pixel_data[47][126] = 0;
        pixel_data[47][127] = 0;
        pixel_data[47][128] = 0;
        pixel_data[47][129] = 0;
        pixel_data[47][130] = 0;
        pixel_data[47][131] = 0;
        pixel_data[47][132] = 0;
        pixel_data[47][133] = 0;
        pixel_data[47][134] = 0;
        pixel_data[47][135] = 0;
        pixel_data[47][136] = 0;
        pixel_data[47][137] = 0;
        pixel_data[47][138] = 0;
        pixel_data[47][139] = 0;
        pixel_data[47][140] = 0;
        pixel_data[47][141] = 0;
        pixel_data[47][142] = 0;
        pixel_data[47][143] = 0;
        pixel_data[47][144] = 0;
        pixel_data[47][145] = 0;
        pixel_data[47][146] = 0;
        pixel_data[47][147] = 0;
        pixel_data[47][148] = 0;
        pixel_data[47][149] = 0;
        pixel_data[47][150] = 0;
        pixel_data[47][151] = 0;
        pixel_data[47][152] = 0;
        pixel_data[47][153] = 0;
        pixel_data[47][154] = 0;
        pixel_data[47][155] = 0;
        pixel_data[47][156] = 0;
        pixel_data[47][157] = 0;
        pixel_data[47][158] = 0;
        pixel_data[47][159] = 0;
        pixel_data[47][160] = 0;
        pixel_data[47][161] = 0;
        pixel_data[47][162] = 0;
        pixel_data[47][163] = 0;
        pixel_data[47][164] = 0;
        pixel_data[47][165] = 0;
        pixel_data[47][166] = 0;
        pixel_data[47][167] = 0;
        pixel_data[47][168] = 0;
        pixel_data[47][169] = 0;
        pixel_data[47][170] = 0;
        pixel_data[47][171] = 0;
        pixel_data[47][172] = 0;
        pixel_data[47][173] = 0;
        pixel_data[47][174] = 0;
        pixel_data[47][175] = 0;
        pixel_data[47][176] = 0;
        pixel_data[47][177] = 0;
        pixel_data[47][178] = 0;
        pixel_data[47][179] = 0;
        pixel_data[47][180] = 0;
        pixel_data[47][181] = 0;
        pixel_data[47][182] = 0;
        pixel_data[47][183] = 0;
        pixel_data[47][184] = 0;
        pixel_data[47][185] = 0;
        pixel_data[47][186] = 0;
        pixel_data[47][187] = 0;
        pixel_data[47][188] = 0;
        pixel_data[47][189] = 0;
        pixel_data[47][190] = 0;
        pixel_data[47][191] = 0;
        pixel_data[47][192] = 0;
        pixel_data[47][193] = 0;
        pixel_data[47][194] = 0;
        pixel_data[47][195] = 0;
        pixel_data[47][196] = 0;
        pixel_data[47][197] = 0;
        pixel_data[47][198] = 0;
        pixel_data[47][199] = 0; // y=47
        pixel_data[48][0] = 0;
        pixel_data[48][1] = 0;
        pixel_data[48][2] = 0;
        pixel_data[48][3] = 0;
        pixel_data[48][4] = 0;
        pixel_data[48][5] = 0;
        pixel_data[48][6] = 0;
        pixel_data[48][7] = 0;
        pixel_data[48][8] = 0;
        pixel_data[48][9] = 0;
        pixel_data[48][10] = 0;
        pixel_data[48][11] = 0;
        pixel_data[48][12] = 0;
        pixel_data[48][13] = 0;
        pixel_data[48][14] = 0;
        pixel_data[48][15] = 0;
        pixel_data[48][16] = 0;
        pixel_data[48][17] = 0;
        pixel_data[48][18] = 0;
        pixel_data[48][19] = 0;
        pixel_data[48][20] = 0;
        pixel_data[48][21] = 0;
        pixel_data[48][22] = 0;
        pixel_data[48][23] = 0;
        pixel_data[48][24] = 0;
        pixel_data[48][25] = 0;
        pixel_data[48][26] = 0;
        pixel_data[48][27] = 0;
        pixel_data[48][28] = 0;
        pixel_data[48][29] = 0;
        pixel_data[48][30] = 0;
        pixel_data[48][31] = 0;
        pixel_data[48][32] = 0;
        pixel_data[48][33] = 0;
        pixel_data[48][34] = 0;
        pixel_data[48][35] = 0;
        pixel_data[48][36] = 0;
        pixel_data[48][37] = 0;
        pixel_data[48][38] = 0;
        pixel_data[48][39] = 0;
        pixel_data[48][40] = 0;
        pixel_data[48][41] = 0;
        pixel_data[48][42] = 0;
        pixel_data[48][43] = 0;
        pixel_data[48][44] = 0;
        pixel_data[48][45] = 0;
        pixel_data[48][46] = 0;
        pixel_data[48][47] = 0;
        pixel_data[48][48] = 0;
        pixel_data[48][49] = 0;
        pixel_data[48][50] = 0;
        pixel_data[48][51] = 0;
        pixel_data[48][52] = 0;
        pixel_data[48][53] = 0;
        pixel_data[48][54] = 0;
        pixel_data[48][55] = 0;
        pixel_data[48][56] = 0;
        pixel_data[48][57] = 0;
        pixel_data[48][58] = 0;
        pixel_data[48][59] = 0;
        pixel_data[48][60] = 0;
        pixel_data[48][61] = 0;
        pixel_data[48][62] = 0;
        pixel_data[48][63] = 0;
        pixel_data[48][64] = 0;
        pixel_data[48][65] = 0;
        pixel_data[48][66] = 0;
        pixel_data[48][67] = 0;
        pixel_data[48][68] = 0;
        pixel_data[48][69] = 0;
        pixel_data[48][70] = 0;
        pixel_data[48][71] = 0;
        pixel_data[48][72] = 0;
        pixel_data[48][73] = 0;
        pixel_data[48][74] = 0;
        pixel_data[48][75] = 0;
        pixel_data[48][76] = 0;
        pixel_data[48][77] = 0;
        pixel_data[48][78] = 0;
        pixel_data[48][79] = 0;
        pixel_data[48][80] = 0;
        pixel_data[48][81] = 0;
        pixel_data[48][82] = 0;
        pixel_data[48][83] = 0;
        pixel_data[48][84] = 0;
        pixel_data[48][85] = 0;
        pixel_data[48][86] = 0;
        pixel_data[48][87] = 0;
        pixel_data[48][88] = 0;
        pixel_data[48][89] = 0;
        pixel_data[48][90] = 0;
        pixel_data[48][91] = 0;
        pixel_data[48][92] = 0;
        pixel_data[48][93] = 0;
        pixel_data[48][94] = 0;
        pixel_data[48][95] = 0;
        pixel_data[48][96] = 0;
        pixel_data[48][97] = 0;
        pixel_data[48][98] = 0;
        pixel_data[48][99] = 0;
        pixel_data[48][100] = 0;
        pixel_data[48][101] = 0;
        pixel_data[48][102] = 0;
        pixel_data[48][103] = 0;
        pixel_data[48][104] = 0;
        pixel_data[48][105] = 0;
        pixel_data[48][106] = 0;
        pixel_data[48][107] = 0;
        pixel_data[48][108] = 0;
        pixel_data[48][109] = 0;
        pixel_data[48][110] = 0;
        pixel_data[48][111] = 0;
        pixel_data[48][112] = 0;
        pixel_data[48][113] = 0;
        pixel_data[48][114] = 0;
        pixel_data[48][115] = 0;
        pixel_data[48][116] = 0;
        pixel_data[48][117] = 0;
        pixel_data[48][118] = 0;
        pixel_data[48][119] = 0;
        pixel_data[48][120] = 0;
        pixel_data[48][121] = 0;
        pixel_data[48][122] = 0;
        pixel_data[48][123] = 0;
        pixel_data[48][124] = 0;
        pixel_data[48][125] = 0;
        pixel_data[48][126] = 0;
        pixel_data[48][127] = 0;
        pixel_data[48][128] = 0;
        pixel_data[48][129] = 0;
        pixel_data[48][130] = 0;
        pixel_data[48][131] = 0;
        pixel_data[48][132] = 0;
        pixel_data[48][133] = 0;
        pixel_data[48][134] = 0;
        pixel_data[48][135] = 0;
        pixel_data[48][136] = 0;
        pixel_data[48][137] = 0;
        pixel_data[48][138] = 0;
        pixel_data[48][139] = 0;
        pixel_data[48][140] = 0;
        pixel_data[48][141] = 0;
        pixel_data[48][142] = 0;
        pixel_data[48][143] = 0;
        pixel_data[48][144] = 0;
        pixel_data[48][145] = 0;
        pixel_data[48][146] = 0;
        pixel_data[48][147] = 0;
        pixel_data[48][148] = 0;
        pixel_data[48][149] = 0;
        pixel_data[48][150] = 0;
        pixel_data[48][151] = 0;
        pixel_data[48][152] = 0;
        pixel_data[48][153] = 0;
        pixel_data[48][154] = 0;
        pixel_data[48][155] = 0;
        pixel_data[48][156] = 0;
        pixel_data[48][157] = 0;
        pixel_data[48][158] = 0;
        pixel_data[48][159] = 0;
        pixel_data[48][160] = 0;
        pixel_data[48][161] = 0;
        pixel_data[48][162] = 0;
        pixel_data[48][163] = 0;
        pixel_data[48][164] = 0;
        pixel_data[48][165] = 0;
        pixel_data[48][166] = 0;
        pixel_data[48][167] = 0;
        pixel_data[48][168] = 0;
        pixel_data[48][169] = 0;
        pixel_data[48][170] = 0;
        pixel_data[48][171] = 0;
        pixel_data[48][172] = 0;
        pixel_data[48][173] = 0;
        pixel_data[48][174] = 0;
        pixel_data[48][175] = 0;
        pixel_data[48][176] = 0;
        pixel_data[48][177] = 0;
        pixel_data[48][178] = 0;
        pixel_data[48][179] = 0;
        pixel_data[48][180] = 0;
        pixel_data[48][181] = 0;
        pixel_data[48][182] = 0;
        pixel_data[48][183] = 0;
        pixel_data[48][184] = 0;
        pixel_data[48][185] = 0;
        pixel_data[48][186] = 0;
        pixel_data[48][187] = 0;
        pixel_data[48][188] = 0;
        pixel_data[48][189] = 0;
        pixel_data[48][190] = 0;
        pixel_data[48][191] = 0;
        pixel_data[48][192] = 0;
        pixel_data[48][193] = 0;
        pixel_data[48][194] = 0;
        pixel_data[48][195] = 0;
        pixel_data[48][196] = 0;
        pixel_data[48][197] = 0;
        pixel_data[48][198] = 0;
        pixel_data[48][199] = 0; // y=48
        pixel_data[49][0] = 0;
        pixel_data[49][1] = 0;
        pixel_data[49][2] = 0;
        pixel_data[49][3] = 0;
        pixel_data[49][4] = 0;
        pixel_data[49][5] = 0;
        pixel_data[49][6] = 0;
        pixel_data[49][7] = 0;
        pixel_data[49][8] = 0;
        pixel_data[49][9] = 0;
        pixel_data[49][10] = 0;
        pixel_data[49][11] = 0;
        pixel_data[49][12] = 0;
        pixel_data[49][13] = 0;
        pixel_data[49][14] = 0;
        pixel_data[49][15] = 0;
        pixel_data[49][16] = 0;
        pixel_data[49][17] = 0;
        pixel_data[49][18] = 0;
        pixel_data[49][19] = 0;
        pixel_data[49][20] = 0;
        pixel_data[49][21] = 0;
        pixel_data[49][22] = 0;
        pixel_data[49][23] = 0;
        pixel_data[49][24] = 0;
        pixel_data[49][25] = 0;
        pixel_data[49][26] = 0;
        pixel_data[49][27] = 0;
        pixel_data[49][28] = 0;
        pixel_data[49][29] = 0;
        pixel_data[49][30] = 0;
        pixel_data[49][31] = 0;
        pixel_data[49][32] = 0;
        pixel_data[49][33] = 0;
        pixel_data[49][34] = 0;
        pixel_data[49][35] = 0;
        pixel_data[49][36] = 0;
        pixel_data[49][37] = 0;
        pixel_data[49][38] = 0;
        pixel_data[49][39] = 0;
        pixel_data[49][40] = 0;
        pixel_data[49][41] = 0;
        pixel_data[49][42] = 0;
        pixel_data[49][43] = 0;
        pixel_data[49][44] = 0;
        pixel_data[49][45] = 0;
        pixel_data[49][46] = 0;
        pixel_data[49][47] = 0;
        pixel_data[49][48] = 0;
        pixel_data[49][49] = 0;
        pixel_data[49][50] = 0;
        pixel_data[49][51] = 0;
        pixel_data[49][52] = 0;
        pixel_data[49][53] = 0;
        pixel_data[49][54] = 0;
        pixel_data[49][55] = 0;
        pixel_data[49][56] = 0;
        pixel_data[49][57] = 0;
        pixel_data[49][58] = 0;
        pixel_data[49][59] = 0;
        pixel_data[49][60] = 0;
        pixel_data[49][61] = 0;
        pixel_data[49][62] = 0;
        pixel_data[49][63] = 0;
        pixel_data[49][64] = 0;
        pixel_data[49][65] = 0;
        pixel_data[49][66] = 0;
        pixel_data[49][67] = 0;
        pixel_data[49][68] = 0;
        pixel_data[49][69] = 0;
        pixel_data[49][70] = 0;
        pixel_data[49][71] = 0;
        pixel_data[49][72] = 0;
        pixel_data[49][73] = 0;
        pixel_data[49][74] = 0;
        pixel_data[49][75] = 0;
        pixel_data[49][76] = 0;
        pixel_data[49][77] = 0;
        pixel_data[49][78] = 0;
        pixel_data[49][79] = 0;
        pixel_data[49][80] = 0;
        pixel_data[49][81] = 0;
        pixel_data[49][82] = 0;
        pixel_data[49][83] = 0;
        pixel_data[49][84] = 0;
        pixel_data[49][85] = 0;
        pixel_data[49][86] = 0;
        pixel_data[49][87] = 0;
        pixel_data[49][88] = 0;
        pixel_data[49][89] = 0;
        pixel_data[49][90] = 0;
        pixel_data[49][91] = 0;
        pixel_data[49][92] = 0;
        pixel_data[49][93] = 0;
        pixel_data[49][94] = 0;
        pixel_data[49][95] = 0;
        pixel_data[49][96] = 0;
        pixel_data[49][97] = 0;
        pixel_data[49][98] = 0;
        pixel_data[49][99] = 0;
        pixel_data[49][100] = 0;
        pixel_data[49][101] = 0;
        pixel_data[49][102] = 0;
        pixel_data[49][103] = 0;
        pixel_data[49][104] = 0;
        pixel_data[49][105] = 0;
        pixel_data[49][106] = 0;
        pixel_data[49][107] = 0;
        pixel_data[49][108] = 0;
        pixel_data[49][109] = 0;
        pixel_data[49][110] = 0;
        pixel_data[49][111] = 0;
        pixel_data[49][112] = 0;
        pixel_data[49][113] = 0;
        pixel_data[49][114] = 0;
        pixel_data[49][115] = 0;
        pixel_data[49][116] = 0;
        pixel_data[49][117] = 0;
        pixel_data[49][118] = 0;
        pixel_data[49][119] = 0;
        pixel_data[49][120] = 0;
        pixel_data[49][121] = 0;
        pixel_data[49][122] = 0;
        pixel_data[49][123] = 0;
        pixel_data[49][124] = 0;
        pixel_data[49][125] = 0;
        pixel_data[49][126] = 0;
        pixel_data[49][127] = 0;
        pixel_data[49][128] = 0;
        pixel_data[49][129] = 0;
        pixel_data[49][130] = 0;
        pixel_data[49][131] = 0;
        pixel_data[49][132] = 0;
        pixel_data[49][133] = 0;
        pixel_data[49][134] = 0;
        pixel_data[49][135] = 0;
        pixel_data[49][136] = 0;
        pixel_data[49][137] = 0;
        pixel_data[49][138] = 0;
        pixel_data[49][139] = 0;
        pixel_data[49][140] = 0;
        pixel_data[49][141] = 0;
        pixel_data[49][142] = 0;
        pixel_data[49][143] = 0;
        pixel_data[49][144] = 0;
        pixel_data[49][145] = 0;
        pixel_data[49][146] = 0;
        pixel_data[49][147] = 0;
        pixel_data[49][148] = 0;
        pixel_data[49][149] = 0;
        pixel_data[49][150] = 0;
        pixel_data[49][151] = 0;
        pixel_data[49][152] = 0;
        pixel_data[49][153] = 0;
        pixel_data[49][154] = 0;
        pixel_data[49][155] = 0;
        pixel_data[49][156] = 0;
        pixel_data[49][157] = 0;
        pixel_data[49][158] = 0;
        pixel_data[49][159] = 0;
        pixel_data[49][160] = 0;
        pixel_data[49][161] = 0;
        pixel_data[49][162] = 0;
        pixel_data[49][163] = 0;
        pixel_data[49][164] = 0;
        pixel_data[49][165] = 0;
        pixel_data[49][166] = 0;
        pixel_data[49][167] = 0;
        pixel_data[49][168] = 0;
        pixel_data[49][169] = 0;
        pixel_data[49][170] = 0;
        pixel_data[49][171] = 0;
        pixel_data[49][172] = 0;
        pixel_data[49][173] = 0;
        pixel_data[49][174] = 0;
        pixel_data[49][175] = 0;
        pixel_data[49][176] = 0;
        pixel_data[49][177] = 0;
        pixel_data[49][178] = 0;
        pixel_data[49][179] = 0;
        pixel_data[49][180] = 0;
        pixel_data[49][181] = 0;
        pixel_data[49][182] = 0;
        pixel_data[49][183] = 0;
        pixel_data[49][184] = 0;
        pixel_data[49][185] = 0;
        pixel_data[49][186] = 0;
        pixel_data[49][187] = 0;
        pixel_data[49][188] = 0;
        pixel_data[49][189] = 0;
        pixel_data[49][190] = 0;
        pixel_data[49][191] = 0;
        pixel_data[49][192] = 0;
        pixel_data[49][193] = 0;
        pixel_data[49][194] = 0;
        pixel_data[49][195] = 0;
        pixel_data[49][196] = 0;
        pixel_data[49][197] = 0;
        pixel_data[49][198] = 0;
        pixel_data[49][199] = 0; // y=49
        pixel_data[50][0] = 0;
        pixel_data[50][1] = 0;
        pixel_data[50][2] = 0;
        pixel_data[50][3] = 0;
        pixel_data[50][4] = 0;
        pixel_data[50][5] = 0;
        pixel_data[50][6] = 0;
        pixel_data[50][7] = 0;
        pixel_data[50][8] = 0;
        pixel_data[50][9] = 0;
        pixel_data[50][10] = 0;
        pixel_data[50][11] = 0;
        pixel_data[50][12] = 0;
        pixel_data[50][13] = 0;
        pixel_data[50][14] = 0;
        pixel_data[50][15] = 0;
        pixel_data[50][16] = 0;
        pixel_data[50][17] = 0;
        pixel_data[50][18] = 0;
        pixel_data[50][19] = 0;
        pixel_data[50][20] = 0;
        pixel_data[50][21] = 0;
        pixel_data[50][22] = 0;
        pixel_data[50][23] = 0;
        pixel_data[50][24] = 0;
        pixel_data[50][25] = 0;
        pixel_data[50][26] = 0;
        pixel_data[50][27] = 0;
        pixel_data[50][28] = 0;
        pixel_data[50][29] = 0;
        pixel_data[50][30] = 0;
        pixel_data[50][31] = 0;
        pixel_data[50][32] = 0;
        pixel_data[50][33] = 0;
        pixel_data[50][34] = 0;
        pixel_data[50][35] = 0;
        pixel_data[50][36] = 0;
        pixel_data[50][37] = 0;
        pixel_data[50][38] = 0;
        pixel_data[50][39] = 0;
        pixel_data[50][40] = 0;
        pixel_data[50][41] = 0;
        pixel_data[50][42] = 0;
        pixel_data[50][43] = 0;
        pixel_data[50][44] = 0;
        pixel_data[50][45] = 0;
        pixel_data[50][46] = 0;
        pixel_data[50][47] = 0;
        pixel_data[50][48] = 0;
        pixel_data[50][49] = 0;
        pixel_data[50][50] = 0;
        pixel_data[50][51] = 0;
        pixel_data[50][52] = 0;
        pixel_data[50][53] = 0;
        pixel_data[50][54] = 0;
        pixel_data[50][55] = 0;
        pixel_data[50][56] = 0;
        pixel_data[50][57] = 0;
        pixel_data[50][58] = 0;
        pixel_data[50][59] = 0;
        pixel_data[50][60] = 0;
        pixel_data[50][61] = 0;
        pixel_data[50][62] = 0;
        pixel_data[50][63] = 0;
        pixel_data[50][64] = 0;
        pixel_data[50][65] = 0;
        pixel_data[50][66] = 0;
        pixel_data[50][67] = 0;
        pixel_data[50][68] = 0;
        pixel_data[50][69] = 0;
        pixel_data[50][70] = 0;
        pixel_data[50][71] = 0;
        pixel_data[50][72] = 0;
        pixel_data[50][73] = 0;
        pixel_data[50][74] = 0;
        pixel_data[50][75] = 0;
        pixel_data[50][76] = 0;
        pixel_data[50][77] = 0;
        pixel_data[50][78] = 0;
        pixel_data[50][79] = 0;
        pixel_data[50][80] = 0;
        pixel_data[50][81] = 0;
        pixel_data[50][82] = 0;
        pixel_data[50][83] = 0;
        pixel_data[50][84] = 0;
        pixel_data[50][85] = 0;
        pixel_data[50][86] = 0;
        pixel_data[50][87] = 0;
        pixel_data[50][88] = 0;
        pixel_data[50][89] = 0;
        pixel_data[50][90] = 0;
        pixel_data[50][91] = 0;
        pixel_data[50][92] = 0;
        pixel_data[50][93] = 0;
        pixel_data[50][94] = 0;
        pixel_data[50][95] = 0;
        pixel_data[50][96] = 0;
        pixel_data[50][97] = 0;
        pixel_data[50][98] = 0;
        pixel_data[50][99] = 0;
        pixel_data[50][100] = 0;
        pixel_data[50][101] = 0;
        pixel_data[50][102] = 0;
        pixel_data[50][103] = 0;
        pixel_data[50][104] = 0;
        pixel_data[50][105] = 0;
        pixel_data[50][106] = 0;
        pixel_data[50][107] = 0;
        pixel_data[50][108] = 0;
        pixel_data[50][109] = 0;
        pixel_data[50][110] = 0;
        pixel_data[50][111] = 0;
        pixel_data[50][112] = 0;
        pixel_data[50][113] = 0;
        pixel_data[50][114] = 0;
        pixel_data[50][115] = 0;
        pixel_data[50][116] = 0;
        pixel_data[50][117] = 0;
        pixel_data[50][118] = 0;
        pixel_data[50][119] = 0;
        pixel_data[50][120] = 0;
        pixel_data[50][121] = 0;
        pixel_data[50][122] = 0;
        pixel_data[50][123] = 0;
        pixel_data[50][124] = 0;
        pixel_data[50][125] = 0;
        pixel_data[50][126] = 0;
        pixel_data[50][127] = 0;
        pixel_data[50][128] = 0;
        pixel_data[50][129] = 0;
        pixel_data[50][130] = 0;
        pixel_data[50][131] = 0;
        pixel_data[50][132] = 0;
        pixel_data[50][133] = 0;
        pixel_data[50][134] = 0;
        pixel_data[50][135] = 0;
        pixel_data[50][136] = 0;
        pixel_data[50][137] = 0;
        pixel_data[50][138] = 0;
        pixel_data[50][139] = 0;
        pixel_data[50][140] = 0;
        pixel_data[50][141] = 0;
        pixel_data[50][142] = 0;
        pixel_data[50][143] = 0;
        pixel_data[50][144] = 0;
        pixel_data[50][145] = 0;
        pixel_data[50][146] = 0;
        pixel_data[50][147] = 0;
        pixel_data[50][148] = 0;
        pixel_data[50][149] = 0;
        pixel_data[50][150] = 0;
        pixel_data[50][151] = 0;
        pixel_data[50][152] = 0;
        pixel_data[50][153] = 0;
        pixel_data[50][154] = 0;
        pixel_data[50][155] = 0;
        pixel_data[50][156] = 0;
        pixel_data[50][157] = 0;
        pixel_data[50][158] = 0;
        pixel_data[50][159] = 0;
        pixel_data[50][160] = 0;
        pixel_data[50][161] = 0;
        pixel_data[50][162] = 0;
        pixel_data[50][163] = 0;
        pixel_data[50][164] = 0;
        pixel_data[50][165] = 0;
        pixel_data[50][166] = 0;
        pixel_data[50][167] = 0;
        pixel_data[50][168] = 0;
        pixel_data[50][169] = 0;
        pixel_data[50][170] = 0;
        pixel_data[50][171] = 0;
        pixel_data[50][172] = 0;
        pixel_data[50][173] = 0;
        pixel_data[50][174] = 0;
        pixel_data[50][175] = 0;
        pixel_data[50][176] = 0;
        pixel_data[50][177] = 0;
        pixel_data[50][178] = 0;
        pixel_data[50][179] = 0;
        pixel_data[50][180] = 0;
        pixel_data[50][181] = 0;
        pixel_data[50][182] = 0;
        pixel_data[50][183] = 0;
        pixel_data[50][184] = 0;
        pixel_data[50][185] = 0;
        pixel_data[50][186] = 0;
        pixel_data[50][187] = 0;
        pixel_data[50][188] = 0;
        pixel_data[50][189] = 0;
        pixel_data[50][190] = 0;
        pixel_data[50][191] = 0;
        pixel_data[50][192] = 0;
        pixel_data[50][193] = 0;
        pixel_data[50][194] = 0;
        pixel_data[50][195] = 0;
        pixel_data[50][196] = 0;
        pixel_data[50][197] = 0;
        pixel_data[50][198] = 0;
        pixel_data[50][199] = 0; // y=50
        pixel_data[51][0] = 0;
        pixel_data[51][1] = 0;
        pixel_data[51][2] = 0;
        pixel_data[51][3] = 0;
        pixel_data[51][4] = 0;
        pixel_data[51][5] = 0;
        pixel_data[51][6] = 0;
        pixel_data[51][7] = 0;
        pixel_data[51][8] = 0;
        pixel_data[51][9] = 0;
        pixel_data[51][10] = 0;
        pixel_data[51][11] = 0;
        pixel_data[51][12] = 0;
        pixel_data[51][13] = 0;
        pixel_data[51][14] = 0;
        pixel_data[51][15] = 0;
        pixel_data[51][16] = 0;
        pixel_data[51][17] = 0;
        pixel_data[51][18] = 0;
        pixel_data[51][19] = 0;
        pixel_data[51][20] = 0;
        pixel_data[51][21] = 0;
        pixel_data[51][22] = 0;
        pixel_data[51][23] = 0;
        pixel_data[51][24] = 0;
        pixel_data[51][25] = 0;
        pixel_data[51][26] = 0;
        pixel_data[51][27] = 0;
        pixel_data[51][28] = 0;
        pixel_data[51][29] = 0;
        pixel_data[51][30] = 0;
        pixel_data[51][31] = 0;
        pixel_data[51][32] = 0;
        pixel_data[51][33] = 0;
        pixel_data[51][34] = 0;
        pixel_data[51][35] = 0;
        pixel_data[51][36] = 0;
        pixel_data[51][37] = 0;
        pixel_data[51][38] = 0;
        pixel_data[51][39] = 0;
        pixel_data[51][40] = 0;
        pixel_data[51][41] = 0;
        pixel_data[51][42] = 0;
        pixel_data[51][43] = 0;
        pixel_data[51][44] = 0;
        pixel_data[51][45] = 0;
        pixel_data[51][46] = 0;
        pixel_data[51][47] = 0;
        pixel_data[51][48] = 0;
        pixel_data[51][49] = 0;
        pixel_data[51][50] = 0;
        pixel_data[51][51] = 0;
        pixel_data[51][52] = 0;
        pixel_data[51][53] = 0;
        pixel_data[51][54] = 0;
        pixel_data[51][55] = 0;
        pixel_data[51][56] = 0;
        pixel_data[51][57] = 0;
        pixel_data[51][58] = 0;
        pixel_data[51][59] = 0;
        pixel_data[51][60] = 0;
        pixel_data[51][61] = 0;
        pixel_data[51][62] = 0;
        pixel_data[51][63] = 0;
        pixel_data[51][64] = 0;
        pixel_data[51][65] = 0;
        pixel_data[51][66] = 0;
        pixel_data[51][67] = 0;
        pixel_data[51][68] = 0;
        pixel_data[51][69] = 0;
        pixel_data[51][70] = 0;
        pixel_data[51][71] = 0;
        pixel_data[51][72] = 0;
        pixel_data[51][73] = 0;
        pixel_data[51][74] = 0;
        pixel_data[51][75] = 0;
        pixel_data[51][76] = 0;
        pixel_data[51][77] = 0;
        pixel_data[51][78] = 0;
        pixel_data[51][79] = 0;
        pixel_data[51][80] = 0;
        pixel_data[51][81] = 0;
        pixel_data[51][82] = 0;
        pixel_data[51][83] = 0;
        pixel_data[51][84] = 0;
        pixel_data[51][85] = 0;
        pixel_data[51][86] = 0;
        pixel_data[51][87] = 0;
        pixel_data[51][88] = 0;
        pixel_data[51][89] = 0;
        pixel_data[51][90] = 0;
        pixel_data[51][91] = 0;
        pixel_data[51][92] = 0;
        pixel_data[51][93] = 0;
        pixel_data[51][94] = 0;
        pixel_data[51][95] = 0;
        pixel_data[51][96] = 0;
        pixel_data[51][97] = 0;
        pixel_data[51][98] = 0;
        pixel_data[51][99] = 0;
        pixel_data[51][100] = 0;
        pixel_data[51][101] = 0;
        pixel_data[51][102] = 0;
        pixel_data[51][103] = 0;
        pixel_data[51][104] = 0;
        pixel_data[51][105] = 0;
        pixel_data[51][106] = 0;
        pixel_data[51][107] = 0;
        pixel_data[51][108] = 0;
        pixel_data[51][109] = 0;
        pixel_data[51][110] = 0;
        pixel_data[51][111] = 0;
        pixel_data[51][112] = 0;
        pixel_data[51][113] = 0;
        pixel_data[51][114] = 0;
        pixel_data[51][115] = 0;
        pixel_data[51][116] = 0;
        pixel_data[51][117] = 0;
        pixel_data[51][118] = 0;
        pixel_data[51][119] = 0;
        pixel_data[51][120] = 0;
        pixel_data[51][121] = 0;
        pixel_data[51][122] = 0;
        pixel_data[51][123] = 0;
        pixel_data[51][124] = 0;
        pixel_data[51][125] = 0;
        pixel_data[51][126] = 0;
        pixel_data[51][127] = 0;
        pixel_data[51][128] = 0;
        pixel_data[51][129] = 0;
        pixel_data[51][130] = 0;
        pixel_data[51][131] = 0;
        pixel_data[51][132] = 0;
        pixel_data[51][133] = 0;
        pixel_data[51][134] = 0;
        pixel_data[51][135] = 0;
        pixel_data[51][136] = 0;
        pixel_data[51][137] = 0;
        pixel_data[51][138] = 0;
        pixel_data[51][139] = 0;
        pixel_data[51][140] = 0;
        pixel_data[51][141] = 0;
        pixel_data[51][142] = 0;
        pixel_data[51][143] = 0;
        pixel_data[51][144] = 0;
        pixel_data[51][145] = 0;
        pixel_data[51][146] = 0;
        pixel_data[51][147] = 0;
        pixel_data[51][148] = 0;
        pixel_data[51][149] = 0;
        pixel_data[51][150] = 0;
        pixel_data[51][151] = 0;
        pixel_data[51][152] = 0;
        pixel_data[51][153] = 0;
        pixel_data[51][154] = 0;
        pixel_data[51][155] = 0;
        pixel_data[51][156] = 0;
        pixel_data[51][157] = 0;
        pixel_data[51][158] = 0;
        pixel_data[51][159] = 0;
        pixel_data[51][160] = 0;
        pixel_data[51][161] = 0;
        pixel_data[51][162] = 0;
        pixel_data[51][163] = 0;
        pixel_data[51][164] = 0;
        pixel_data[51][165] = 0;
        pixel_data[51][166] = 0;
        pixel_data[51][167] = 0;
        pixel_data[51][168] = 0;
        pixel_data[51][169] = 0;
        pixel_data[51][170] = 0;
        pixel_data[51][171] = 0;
        pixel_data[51][172] = 0;
        pixel_data[51][173] = 0;
        pixel_data[51][174] = 0;
        pixel_data[51][175] = 0;
        pixel_data[51][176] = 0;
        pixel_data[51][177] = 0;
        pixel_data[51][178] = 0;
        pixel_data[51][179] = 0;
        pixel_data[51][180] = 0;
        pixel_data[51][181] = 0;
        pixel_data[51][182] = 0;
        pixel_data[51][183] = 0;
        pixel_data[51][184] = 0;
        pixel_data[51][185] = 0;
        pixel_data[51][186] = 0;
        pixel_data[51][187] = 0;
        pixel_data[51][188] = 0;
        pixel_data[51][189] = 0;
        pixel_data[51][190] = 0;
        pixel_data[51][191] = 0;
        pixel_data[51][192] = 0;
        pixel_data[51][193] = 0;
        pixel_data[51][194] = 0;
        pixel_data[51][195] = 0;
        pixel_data[51][196] = 0;
        pixel_data[51][197] = 0;
        pixel_data[51][198] = 0;
        pixel_data[51][199] = 0; // y=51
        pixel_data[52][0] = 0;
        pixel_data[52][1] = 0;
        pixel_data[52][2] = 0;
        pixel_data[52][3] = 0;
        pixel_data[52][4] = 0;
        pixel_data[52][5] = 0;
        pixel_data[52][6] = 0;
        pixel_data[52][7] = 0;
        pixel_data[52][8] = 0;
        pixel_data[52][9] = 0;
        pixel_data[52][10] = 0;
        pixel_data[52][11] = 0;
        pixel_data[52][12] = 0;
        pixel_data[52][13] = 0;
        pixel_data[52][14] = 0;
        pixel_data[52][15] = 0;
        pixel_data[52][16] = 0;
        pixel_data[52][17] = 0;
        pixel_data[52][18] = 0;
        pixel_data[52][19] = 0;
        pixel_data[52][20] = 0;
        pixel_data[52][21] = 0;
        pixel_data[52][22] = 0;
        pixel_data[52][23] = 0;
        pixel_data[52][24] = 0;
        pixel_data[52][25] = 0;
        pixel_data[52][26] = 0;
        pixel_data[52][27] = 0;
        pixel_data[52][28] = 0;
        pixel_data[52][29] = 0;
        pixel_data[52][30] = 0;
        pixel_data[52][31] = 0;
        pixel_data[52][32] = 0;
        pixel_data[52][33] = 0;
        pixel_data[52][34] = 0;
        pixel_data[52][35] = 0;
        pixel_data[52][36] = 0;
        pixel_data[52][37] = 0;
        pixel_data[52][38] = 0;
        pixel_data[52][39] = 0;
        pixel_data[52][40] = 0;
        pixel_data[52][41] = 0;
        pixel_data[52][42] = 0;
        pixel_data[52][43] = 0;
        pixel_data[52][44] = 0;
        pixel_data[52][45] = 0;
        pixel_data[52][46] = 0;
        pixel_data[52][47] = 0;
        pixel_data[52][48] = 0;
        pixel_data[52][49] = 0;
        pixel_data[52][50] = 0;
        pixel_data[52][51] = 0;
        pixel_data[52][52] = 0;
        pixel_data[52][53] = 0;
        pixel_data[52][54] = 0;
        pixel_data[52][55] = 0;
        pixel_data[52][56] = 0;
        pixel_data[52][57] = 0;
        pixel_data[52][58] = 0;
        pixel_data[52][59] = 0;
        pixel_data[52][60] = 0;
        pixel_data[52][61] = 0;
        pixel_data[52][62] = 0;
        pixel_data[52][63] = 0;
        pixel_data[52][64] = 0;
        pixel_data[52][65] = 0;
        pixel_data[52][66] = 0;
        pixel_data[52][67] = 0;
        pixel_data[52][68] = 0;
        pixel_data[52][69] = 0;
        pixel_data[52][70] = 0;
        pixel_data[52][71] = 0;
        pixel_data[52][72] = 0;
        pixel_data[52][73] = 0;
        pixel_data[52][74] = 0;
        pixel_data[52][75] = 0;
        pixel_data[52][76] = 0;
        pixel_data[52][77] = 0;
        pixel_data[52][78] = 0;
        pixel_data[52][79] = 0;
        pixel_data[52][80] = 0;
        pixel_data[52][81] = 0;
        pixel_data[52][82] = 0;
        pixel_data[52][83] = 0;
        pixel_data[52][84] = 0;
        pixel_data[52][85] = 0;
        pixel_data[52][86] = 0;
        pixel_data[52][87] = 0;
        pixel_data[52][88] = 0;
        pixel_data[52][89] = 0;
        pixel_data[52][90] = 0;
        pixel_data[52][91] = 0;
        pixel_data[52][92] = 0;
        pixel_data[52][93] = 0;
        pixel_data[52][94] = 0;
        pixel_data[52][95] = 0;
        pixel_data[52][96] = 0;
        pixel_data[52][97] = 0;
        pixel_data[52][98] = 0;
        pixel_data[52][99] = 0;
        pixel_data[52][100] = 0;
        pixel_data[52][101] = 0;
        pixel_data[52][102] = 0;
        pixel_data[52][103] = 0;
        pixel_data[52][104] = 0;
        pixel_data[52][105] = 0;
        pixel_data[52][106] = 0;
        pixel_data[52][107] = 0;
        pixel_data[52][108] = 0;
        pixel_data[52][109] = 0;
        pixel_data[52][110] = 0;
        pixel_data[52][111] = 0;
        pixel_data[52][112] = 0;
        pixel_data[52][113] = 0;
        pixel_data[52][114] = 0;
        pixel_data[52][115] = 0;
        pixel_data[52][116] = 0;
        pixel_data[52][117] = 0;
        pixel_data[52][118] = 0;
        pixel_data[52][119] = 0;
        pixel_data[52][120] = 0;
        pixel_data[52][121] = 0;
        pixel_data[52][122] = 0;
        pixel_data[52][123] = 0;
        pixel_data[52][124] = 0;
        pixel_data[52][125] = 0;
        pixel_data[52][126] = 0;
        pixel_data[52][127] = 0;
        pixel_data[52][128] = 0;
        pixel_data[52][129] = 0;
        pixel_data[52][130] = 0;
        pixel_data[52][131] = 0;
        pixel_data[52][132] = 0;
        pixel_data[52][133] = 0;
        pixel_data[52][134] = 0;
        pixel_data[52][135] = 0;
        pixel_data[52][136] = 0;
        pixel_data[52][137] = 0;
        pixel_data[52][138] = 0;
        pixel_data[52][139] = 0;
        pixel_data[52][140] = 0;
        pixel_data[52][141] = 0;
        pixel_data[52][142] = 0;
        pixel_data[52][143] = 0;
        pixel_data[52][144] = 0;
        pixel_data[52][145] = 0;
        pixel_data[52][146] = 0;
        pixel_data[52][147] = 0;
        pixel_data[52][148] = 0;
        pixel_data[52][149] = 0;
        pixel_data[52][150] = 0;
        pixel_data[52][151] = 0;
        pixel_data[52][152] = 0;
        pixel_data[52][153] = 0;
        pixel_data[52][154] = 0;
        pixel_data[52][155] = 0;
        pixel_data[52][156] = 0;
        pixel_data[52][157] = 0;
        pixel_data[52][158] = 0;
        pixel_data[52][159] = 0;
        pixel_data[52][160] = 0;
        pixel_data[52][161] = 0;
        pixel_data[52][162] = 0;
        pixel_data[52][163] = 0;
        pixel_data[52][164] = 0;
        pixel_data[52][165] = 0;
        pixel_data[52][166] = 0;
        pixel_data[52][167] = 0;
        pixel_data[52][168] = 0;
        pixel_data[52][169] = 0;
        pixel_data[52][170] = 0;
        pixel_data[52][171] = 0;
        pixel_data[52][172] = 0;
        pixel_data[52][173] = 0;
        pixel_data[52][174] = 0;
        pixel_data[52][175] = 0;
        pixel_data[52][176] = 0;
        pixel_data[52][177] = 0;
        pixel_data[52][178] = 0;
        pixel_data[52][179] = 0;
        pixel_data[52][180] = 0;
        pixel_data[52][181] = 0;
        pixel_data[52][182] = 0;
        pixel_data[52][183] = 0;
        pixel_data[52][184] = 0;
        pixel_data[52][185] = 0;
        pixel_data[52][186] = 0;
        pixel_data[52][187] = 0;
        pixel_data[52][188] = 0;
        pixel_data[52][189] = 0;
        pixel_data[52][190] = 0;
        pixel_data[52][191] = 0;
        pixel_data[52][192] = 0;
        pixel_data[52][193] = 0;
        pixel_data[52][194] = 0;
        pixel_data[52][195] = 0;
        pixel_data[52][196] = 0;
        pixel_data[52][197] = 0;
        pixel_data[52][198] = 0;
        pixel_data[52][199] = 0; // y=52
        pixel_data[53][0] = 0;
        pixel_data[53][1] = 0;
        pixel_data[53][2] = 0;
        pixel_data[53][3] = 0;
        pixel_data[53][4] = 0;
        pixel_data[53][5] = 0;
        pixel_data[53][6] = 0;
        pixel_data[53][7] = 0;
        pixel_data[53][8] = 0;
        pixel_data[53][9] = 0;
        pixel_data[53][10] = 0;
        pixel_data[53][11] = 0;
        pixel_data[53][12] = 0;
        pixel_data[53][13] = 0;
        pixel_data[53][14] = 0;
        pixel_data[53][15] = 0;
        pixel_data[53][16] = 0;
        pixel_data[53][17] = 0;
        pixel_data[53][18] = 0;
        pixel_data[53][19] = 0;
        pixel_data[53][20] = 0;
        pixel_data[53][21] = 0;
        pixel_data[53][22] = 0;
        pixel_data[53][23] = 0;
        pixel_data[53][24] = 0;
        pixel_data[53][25] = 0;
        pixel_data[53][26] = 0;
        pixel_data[53][27] = 0;
        pixel_data[53][28] = 0;
        pixel_data[53][29] = 0;
        pixel_data[53][30] = 0;
        pixel_data[53][31] = 0;
        pixel_data[53][32] = 0;
        pixel_data[53][33] = 0;
        pixel_data[53][34] = 0;
        pixel_data[53][35] = 0;
        pixel_data[53][36] = 0;
        pixel_data[53][37] = 0;
        pixel_data[53][38] = 0;
        pixel_data[53][39] = 0;
        pixel_data[53][40] = 0;
        pixel_data[53][41] = 0;
        pixel_data[53][42] = 0;
        pixel_data[53][43] = 0;
        pixel_data[53][44] = 0;
        pixel_data[53][45] = 0;
        pixel_data[53][46] = 0;
        pixel_data[53][47] = 0;
        pixel_data[53][48] = 0;
        pixel_data[53][49] = 0;
        pixel_data[53][50] = 0;
        pixel_data[53][51] = 0;
        pixel_data[53][52] = 0;
        pixel_data[53][53] = 0;
        pixel_data[53][54] = 0;
        pixel_data[53][55] = 0;
        pixel_data[53][56] = 0;
        pixel_data[53][57] = 0;
        pixel_data[53][58] = 0;
        pixel_data[53][59] = 0;
        pixel_data[53][60] = 0;
        pixel_data[53][61] = 0;
        pixel_data[53][62] = 0;
        pixel_data[53][63] = 0;
        pixel_data[53][64] = 0;
        pixel_data[53][65] = 0;
        pixel_data[53][66] = 0;
        pixel_data[53][67] = 0;
        pixel_data[53][68] = 0;
        pixel_data[53][69] = 0;
        pixel_data[53][70] = 0;
        pixel_data[53][71] = 0;
        pixel_data[53][72] = 0;
        pixel_data[53][73] = 0;
        pixel_data[53][74] = 0;
        pixel_data[53][75] = 0;
        pixel_data[53][76] = 0;
        pixel_data[53][77] = 0;
        pixel_data[53][78] = 0;
        pixel_data[53][79] = 0;
        pixel_data[53][80] = 0;
        pixel_data[53][81] = 0;
        pixel_data[53][82] = 0;
        pixel_data[53][83] = 0;
        pixel_data[53][84] = 0;
        pixel_data[53][85] = 0;
        pixel_data[53][86] = 0;
        pixel_data[53][87] = 0;
        pixel_data[53][88] = 0;
        pixel_data[53][89] = 0;
        pixel_data[53][90] = 0;
        pixel_data[53][91] = 0;
        pixel_data[53][92] = 0;
        pixel_data[53][93] = 0;
        pixel_data[53][94] = 0;
        pixel_data[53][95] = 0;
        pixel_data[53][96] = 0;
        pixel_data[53][97] = 0;
        pixel_data[53][98] = 0;
        pixel_data[53][99] = 0;
        pixel_data[53][100] = 0;
        pixel_data[53][101] = 0;
        pixel_data[53][102] = 0;
        pixel_data[53][103] = 0;
        pixel_data[53][104] = 0;
        pixel_data[53][105] = 0;
        pixel_data[53][106] = 0;
        pixel_data[53][107] = 0;
        pixel_data[53][108] = 0;
        pixel_data[53][109] = 0;
        pixel_data[53][110] = 0;
        pixel_data[53][111] = 0;
        pixel_data[53][112] = 0;
        pixel_data[53][113] = 0;
        pixel_data[53][114] = 0;
        pixel_data[53][115] = 0;
        pixel_data[53][116] = 0;
        pixel_data[53][117] = 0;
        pixel_data[53][118] = 0;
        pixel_data[53][119] = 0;
        pixel_data[53][120] = 0;
        pixel_data[53][121] = 0;
        pixel_data[53][122] = 0;
        pixel_data[53][123] = 0;
        pixel_data[53][124] = 0;
        pixel_data[53][125] = 0;
        pixel_data[53][126] = 0;
        pixel_data[53][127] = 0;
        pixel_data[53][128] = 0;
        pixel_data[53][129] = 0;
        pixel_data[53][130] = 0;
        pixel_data[53][131] = 0;
        pixel_data[53][132] = 0;
        pixel_data[53][133] = 0;
        pixel_data[53][134] = 0;
        pixel_data[53][135] = 0;
        pixel_data[53][136] = 0;
        pixel_data[53][137] = 0;
        pixel_data[53][138] = 0;
        pixel_data[53][139] = 0;
        pixel_data[53][140] = 0;
        pixel_data[53][141] = 0;
        pixel_data[53][142] = 0;
        pixel_data[53][143] = 0;
        pixel_data[53][144] = 0;
        pixel_data[53][145] = 0;
        pixel_data[53][146] = 0;
        pixel_data[53][147] = 0;
        pixel_data[53][148] = 0;
        pixel_data[53][149] = 0;
        pixel_data[53][150] = 0;
        pixel_data[53][151] = 0;
        pixel_data[53][152] = 0;
        pixel_data[53][153] = 0;
        pixel_data[53][154] = 0;
        pixel_data[53][155] = 0;
        pixel_data[53][156] = 0;
        pixel_data[53][157] = 0;
        pixel_data[53][158] = 0;
        pixel_data[53][159] = 0;
        pixel_data[53][160] = 0;
        pixel_data[53][161] = 0;
        pixel_data[53][162] = 0;
        pixel_data[53][163] = 0;
        pixel_data[53][164] = 0;
        pixel_data[53][165] = 0;
        pixel_data[53][166] = 0;
        pixel_data[53][167] = 0;
        pixel_data[53][168] = 0;
        pixel_data[53][169] = 0;
        pixel_data[53][170] = 0;
        pixel_data[53][171] = 0;
        pixel_data[53][172] = 0;
        pixel_data[53][173] = 0;
        pixel_data[53][174] = 0;
        pixel_data[53][175] = 0;
        pixel_data[53][176] = 0;
        pixel_data[53][177] = 0;
        pixel_data[53][178] = 0;
        pixel_data[53][179] = 0;
        pixel_data[53][180] = 0;
        pixel_data[53][181] = 0;
        pixel_data[53][182] = 0;
        pixel_data[53][183] = 0;
        pixel_data[53][184] = 0;
        pixel_data[53][185] = 0;
        pixel_data[53][186] = 0;
        pixel_data[53][187] = 0;
        pixel_data[53][188] = 0;
        pixel_data[53][189] = 0;
        pixel_data[53][190] = 0;
        pixel_data[53][191] = 0;
        pixel_data[53][192] = 0;
        pixel_data[53][193] = 0;
        pixel_data[53][194] = 0;
        pixel_data[53][195] = 0;
        pixel_data[53][196] = 0;
        pixel_data[53][197] = 0;
        pixel_data[53][198] = 0;
        pixel_data[53][199] = 0; // y=53
        pixel_data[54][0] = 0;
        pixel_data[54][1] = 0;
        pixel_data[54][2] = 0;
        pixel_data[54][3] = 0;
        pixel_data[54][4] = 0;
        pixel_data[54][5] = 0;
        pixel_data[54][6] = 0;
        pixel_data[54][7] = 0;
        pixel_data[54][8] = 0;
        pixel_data[54][9] = 0;
        pixel_data[54][10] = 0;
        pixel_data[54][11] = 0;
        pixel_data[54][12] = 0;
        pixel_data[54][13] = 0;
        pixel_data[54][14] = 0;
        pixel_data[54][15] = 0;
        pixel_data[54][16] = 0;
        pixel_data[54][17] = 0;
        pixel_data[54][18] = 0;
        pixel_data[54][19] = 0;
        pixel_data[54][20] = 0;
        pixel_data[54][21] = 0;
        pixel_data[54][22] = 0;
        pixel_data[54][23] = 0;
        pixel_data[54][24] = 0;
        pixel_data[54][25] = 0;
        pixel_data[54][26] = 0;
        pixel_data[54][27] = 0;
        pixel_data[54][28] = 0;
        pixel_data[54][29] = 0;
        pixel_data[54][30] = 0;
        pixel_data[54][31] = 0;
        pixel_data[54][32] = 0;
        pixel_data[54][33] = 0;
        pixel_data[54][34] = 0;
        pixel_data[54][35] = 0;
        pixel_data[54][36] = 0;
        pixel_data[54][37] = 0;
        pixel_data[54][38] = 0;
        pixel_data[54][39] = 0;
        pixel_data[54][40] = 0;
        pixel_data[54][41] = 0;
        pixel_data[54][42] = 0;
        pixel_data[54][43] = 0;
        pixel_data[54][44] = 0;
        pixel_data[54][45] = 0;
        pixel_data[54][46] = 0;
        pixel_data[54][47] = 0;
        pixel_data[54][48] = 0;
        pixel_data[54][49] = 0;
        pixel_data[54][50] = 0;
        pixel_data[54][51] = 0;
        pixel_data[54][52] = 0;
        pixel_data[54][53] = 0;
        pixel_data[54][54] = 0;
        pixel_data[54][55] = 0;
        pixel_data[54][56] = 0;
        pixel_data[54][57] = 0;
        pixel_data[54][58] = 0;
        pixel_data[54][59] = 0;
        pixel_data[54][60] = 0;
        pixel_data[54][61] = 0;
        pixel_data[54][62] = 0;
        pixel_data[54][63] = 0;
        pixel_data[54][64] = 0;
        pixel_data[54][65] = 0;
        pixel_data[54][66] = 0;
        pixel_data[54][67] = 0;
        pixel_data[54][68] = 0;
        pixel_data[54][69] = 0;
        pixel_data[54][70] = 0;
        pixel_data[54][71] = 0;
        pixel_data[54][72] = 0;
        pixel_data[54][73] = 0;
        pixel_data[54][74] = 0;
        pixel_data[54][75] = 0;
        pixel_data[54][76] = 0;
        pixel_data[54][77] = 0;
        pixel_data[54][78] = 0;
        pixel_data[54][79] = 0;
        pixel_data[54][80] = 0;
        pixel_data[54][81] = 0;
        pixel_data[54][82] = 0;
        pixel_data[54][83] = 0;
        pixel_data[54][84] = 0;
        pixel_data[54][85] = 0;
        pixel_data[54][86] = 0;
        pixel_data[54][87] = 0;
        pixel_data[54][88] = 0;
        pixel_data[54][89] = 0;
        pixel_data[54][90] = 0;
        pixel_data[54][91] = 0;
        pixel_data[54][92] = 0;
        pixel_data[54][93] = 0;
        pixel_data[54][94] = 0;
        pixel_data[54][95] = 0;
        pixel_data[54][96] = 0;
        pixel_data[54][97] = 0;
        pixel_data[54][98] = 0;
        pixel_data[54][99] = 0;
        pixel_data[54][100] = 0;
        pixel_data[54][101] = 0;
        pixel_data[54][102] = 0;
        pixel_data[54][103] = 0;
        pixel_data[54][104] = 0;
        pixel_data[54][105] = 0;
        pixel_data[54][106] = 0;
        pixel_data[54][107] = 0;
        pixel_data[54][108] = 0;
        pixel_data[54][109] = 0;
        pixel_data[54][110] = 0;
        pixel_data[54][111] = 0;
        pixel_data[54][112] = 0;
        pixel_data[54][113] = 0;
        pixel_data[54][114] = 0;
        pixel_data[54][115] = 0;
        pixel_data[54][116] = 0;
        pixel_data[54][117] = 0;
        pixel_data[54][118] = 0;
        pixel_data[54][119] = 0;
        pixel_data[54][120] = 0;
        pixel_data[54][121] = 0;
        pixel_data[54][122] = 0;
        pixel_data[54][123] = 0;
        pixel_data[54][124] = 0;
        pixel_data[54][125] = 0;
        pixel_data[54][126] = 0;
        pixel_data[54][127] = 0;
        pixel_data[54][128] = 0;
        pixel_data[54][129] = 0;
        pixel_data[54][130] = 0;
        pixel_data[54][131] = 0;
        pixel_data[54][132] = 0;
        pixel_data[54][133] = 0;
        pixel_data[54][134] = 0;
        pixel_data[54][135] = 0;
        pixel_data[54][136] = 0;
        pixel_data[54][137] = 0;
        pixel_data[54][138] = 0;
        pixel_data[54][139] = 0;
        pixel_data[54][140] = 0;
        pixel_data[54][141] = 0;
        pixel_data[54][142] = 0;
        pixel_data[54][143] = 0;
        pixel_data[54][144] = 0;
        pixel_data[54][145] = 0;
        pixel_data[54][146] = 0;
        pixel_data[54][147] = 0;
        pixel_data[54][148] = 0;
        pixel_data[54][149] = 0;
        pixel_data[54][150] = 0;
        pixel_data[54][151] = 0;
        pixel_data[54][152] = 0;
        pixel_data[54][153] = 0;
        pixel_data[54][154] = 0;
        pixel_data[54][155] = 0;
        pixel_data[54][156] = 0;
        pixel_data[54][157] = 0;
        pixel_data[54][158] = 0;
        pixel_data[54][159] = 0;
        pixel_data[54][160] = 0;
        pixel_data[54][161] = 0;
        pixel_data[54][162] = 0;
        pixel_data[54][163] = 0;
        pixel_data[54][164] = 0;
        pixel_data[54][165] = 0;
        pixel_data[54][166] = 0;
        pixel_data[54][167] = 0;
        pixel_data[54][168] = 0;
        pixel_data[54][169] = 0;
        pixel_data[54][170] = 0;
        pixel_data[54][171] = 0;
        pixel_data[54][172] = 0;
        pixel_data[54][173] = 0;
        pixel_data[54][174] = 0;
        pixel_data[54][175] = 0;
        pixel_data[54][176] = 0;
        pixel_data[54][177] = 0;
        pixel_data[54][178] = 0;
        pixel_data[54][179] = 0;
        pixel_data[54][180] = 0;
        pixel_data[54][181] = 0;
        pixel_data[54][182] = 0;
        pixel_data[54][183] = 0;
        pixel_data[54][184] = 0;
        pixel_data[54][185] = 0;
        pixel_data[54][186] = 0;
        pixel_data[54][187] = 0;
        pixel_data[54][188] = 0;
        pixel_data[54][189] = 0;
        pixel_data[54][190] = 0;
        pixel_data[54][191] = 0;
        pixel_data[54][192] = 0;
        pixel_data[54][193] = 0;
        pixel_data[54][194] = 0;
        pixel_data[54][195] = 0;
        pixel_data[54][196] = 0;
        pixel_data[54][197] = 0;
        pixel_data[54][198] = 0;
        pixel_data[54][199] = 0; // y=54
        pixel_data[55][0] = 0;
        pixel_data[55][1] = 0;
        pixel_data[55][2] = 0;
        pixel_data[55][3] = 0;
        pixel_data[55][4] = 0;
        pixel_data[55][5] = 0;
        pixel_data[55][6] = 0;
        pixel_data[55][7] = 0;
        pixel_data[55][8] = 0;
        pixel_data[55][9] = 0;
        pixel_data[55][10] = 0;
        pixel_data[55][11] = 0;
        pixel_data[55][12] = 0;
        pixel_data[55][13] = 0;
        pixel_data[55][14] = 0;
        pixel_data[55][15] = 0;
        pixel_data[55][16] = 0;
        pixel_data[55][17] = 0;
        pixel_data[55][18] = 0;
        pixel_data[55][19] = 0;
        pixel_data[55][20] = 0;
        pixel_data[55][21] = 0;
        pixel_data[55][22] = 0;
        pixel_data[55][23] = 0;
        pixel_data[55][24] = 0;
        pixel_data[55][25] = 0;
        pixel_data[55][26] = 0;
        pixel_data[55][27] = 0;
        pixel_data[55][28] = 0;
        pixel_data[55][29] = 0;
        pixel_data[55][30] = 0;
        pixel_data[55][31] = 0;
        pixel_data[55][32] = 0;
        pixel_data[55][33] = 0;
        pixel_data[55][34] = 0;
        pixel_data[55][35] = 0;
        pixel_data[55][36] = 0;
        pixel_data[55][37] = 0;
        pixel_data[55][38] = 0;
        pixel_data[55][39] = 0;
        pixel_data[55][40] = 0;
        pixel_data[55][41] = 0;
        pixel_data[55][42] = 0;
        pixel_data[55][43] = 0;
        pixel_data[55][44] = 0;
        pixel_data[55][45] = 0;
        pixel_data[55][46] = 0;
        pixel_data[55][47] = 0;
        pixel_data[55][48] = 0;
        pixel_data[55][49] = 0;
        pixel_data[55][50] = 0;
        pixel_data[55][51] = 0;
        pixel_data[55][52] = 0;
        pixel_data[55][53] = 0;
        pixel_data[55][54] = 0;
        pixel_data[55][55] = 0;
        pixel_data[55][56] = 0;
        pixel_data[55][57] = 0;
        pixel_data[55][58] = 0;
        pixel_data[55][59] = 0;
        pixel_data[55][60] = 0;
        pixel_data[55][61] = 0;
        pixel_data[55][62] = 0;
        pixel_data[55][63] = 0;
        pixel_data[55][64] = 0;
        pixel_data[55][65] = 0;
        pixel_data[55][66] = 0;
        pixel_data[55][67] = 0;
        pixel_data[55][68] = 0;
        pixel_data[55][69] = 0;
        pixel_data[55][70] = 0;
        pixel_data[55][71] = 0;
        pixel_data[55][72] = 0;
        pixel_data[55][73] = 0;
        pixel_data[55][74] = 0;
        pixel_data[55][75] = 0;
        pixel_data[55][76] = 0;
        pixel_data[55][77] = 0;
        pixel_data[55][78] = 0;
        pixel_data[55][79] = 0;
        pixel_data[55][80] = 0;
        pixel_data[55][81] = 0;
        pixel_data[55][82] = 0;
        pixel_data[55][83] = 0;
        pixel_data[55][84] = 0;
        pixel_data[55][85] = 0;
        pixel_data[55][86] = 0;
        pixel_data[55][87] = 0;
        pixel_data[55][88] = 0;
        pixel_data[55][89] = 0;
        pixel_data[55][90] = 0;
        pixel_data[55][91] = 0;
        pixel_data[55][92] = 0;
        pixel_data[55][93] = 0;
        pixel_data[55][94] = 0;
        pixel_data[55][95] = 0;
        pixel_data[55][96] = 0;
        pixel_data[55][97] = 0;
        pixel_data[55][98] = 0;
        pixel_data[55][99] = 0;
        pixel_data[55][100] = 0;
        pixel_data[55][101] = 0;
        pixel_data[55][102] = 0;
        pixel_data[55][103] = 0;
        pixel_data[55][104] = 0;
        pixel_data[55][105] = 0;
        pixel_data[55][106] = 0;
        pixel_data[55][107] = 0;
        pixel_data[55][108] = 0;
        pixel_data[55][109] = 0;
        pixel_data[55][110] = 0;
        pixel_data[55][111] = 0;
        pixel_data[55][112] = 0;
        pixel_data[55][113] = 0;
        pixel_data[55][114] = 0;
        pixel_data[55][115] = 0;
        pixel_data[55][116] = 0;
        pixel_data[55][117] = 0;
        pixel_data[55][118] = 0;
        pixel_data[55][119] = 0;
        pixel_data[55][120] = 0;
        pixel_data[55][121] = 0;
        pixel_data[55][122] = 0;
        pixel_data[55][123] = 0;
        pixel_data[55][124] = 0;
        pixel_data[55][125] = 0;
        pixel_data[55][126] = 0;
        pixel_data[55][127] = 0;
        pixel_data[55][128] = 0;
        pixel_data[55][129] = 0;
        pixel_data[55][130] = 0;
        pixel_data[55][131] = 0;
        pixel_data[55][132] = 0;
        pixel_data[55][133] = 0;
        pixel_data[55][134] = 0;
        pixel_data[55][135] = 0;
        pixel_data[55][136] = 0;
        pixel_data[55][137] = 0;
        pixel_data[55][138] = 0;
        pixel_data[55][139] = 0;
        pixel_data[55][140] = 0;
        pixel_data[55][141] = 0;
        pixel_data[55][142] = 0;
        pixel_data[55][143] = 0;
        pixel_data[55][144] = 0;
        pixel_data[55][145] = 0;
        pixel_data[55][146] = 0;
        pixel_data[55][147] = 0;
        pixel_data[55][148] = 0;
        pixel_data[55][149] = 0;
        pixel_data[55][150] = 0;
        pixel_data[55][151] = 0;
        pixel_data[55][152] = 0;
        pixel_data[55][153] = 0;
        pixel_data[55][154] = 0;
        pixel_data[55][155] = 0;
        pixel_data[55][156] = 0;
        pixel_data[55][157] = 0;
        pixel_data[55][158] = 0;
        pixel_data[55][159] = 0;
        pixel_data[55][160] = 0;
        pixel_data[55][161] = 0;
        pixel_data[55][162] = 0;
        pixel_data[55][163] = 0;
        pixel_data[55][164] = 0;
        pixel_data[55][165] = 0;
        pixel_data[55][166] = 0;
        pixel_data[55][167] = 0;
        pixel_data[55][168] = 0;
        pixel_data[55][169] = 0;
        pixel_data[55][170] = 0;
        pixel_data[55][171] = 0;
        pixel_data[55][172] = 0;
        pixel_data[55][173] = 0;
        pixel_data[55][174] = 0;
        pixel_data[55][175] = 0;
        pixel_data[55][176] = 0;
        pixel_data[55][177] = 0;
        pixel_data[55][178] = 0;
        pixel_data[55][179] = 0;
        pixel_data[55][180] = 0;
        pixel_data[55][181] = 0;
        pixel_data[55][182] = 0;
        pixel_data[55][183] = 0;
        pixel_data[55][184] = 0;
        pixel_data[55][185] = 0;
        pixel_data[55][186] = 0;
        pixel_data[55][187] = 0;
        pixel_data[55][188] = 0;
        pixel_data[55][189] = 0;
        pixel_data[55][190] = 0;
        pixel_data[55][191] = 0;
        pixel_data[55][192] = 0;
        pixel_data[55][193] = 0;
        pixel_data[55][194] = 0;
        pixel_data[55][195] = 0;
        pixel_data[55][196] = 0;
        pixel_data[55][197] = 0;
        pixel_data[55][198] = 0;
        pixel_data[55][199] = 0; // y=55
        pixel_data[56][0] = 0;
        pixel_data[56][1] = 0;
        pixel_data[56][2] = 0;
        pixel_data[56][3] = 0;
        pixel_data[56][4] = 0;
        pixel_data[56][5] = 0;
        pixel_data[56][6] = 0;
        pixel_data[56][7] = 0;
        pixel_data[56][8] = 0;
        pixel_data[56][9] = 0;
        pixel_data[56][10] = 0;
        pixel_data[56][11] = 0;
        pixel_data[56][12] = 0;
        pixel_data[56][13] = 0;
        pixel_data[56][14] = 0;
        pixel_data[56][15] = 0;
        pixel_data[56][16] = 0;
        pixel_data[56][17] = 0;
        pixel_data[56][18] = 0;
        pixel_data[56][19] = 0;
        pixel_data[56][20] = 0;
        pixel_data[56][21] = 0;
        pixel_data[56][22] = 0;
        pixel_data[56][23] = 0;
        pixel_data[56][24] = 0;
        pixel_data[56][25] = 0;
        pixel_data[56][26] = 0;
        pixel_data[56][27] = 0;
        pixel_data[56][28] = 0;
        pixel_data[56][29] = 0;
        pixel_data[56][30] = 0;
        pixel_data[56][31] = 0;
        pixel_data[56][32] = 0;
        pixel_data[56][33] = 0;
        pixel_data[56][34] = 0;
        pixel_data[56][35] = 0;
        pixel_data[56][36] = 0;
        pixel_data[56][37] = 0;
        pixel_data[56][38] = 0;
        pixel_data[56][39] = 0;
        pixel_data[56][40] = 0;
        pixel_data[56][41] = 0;
        pixel_data[56][42] = 0;
        pixel_data[56][43] = 0;
        pixel_data[56][44] = 0;
        pixel_data[56][45] = 0;
        pixel_data[56][46] = 0;
        pixel_data[56][47] = 0;
        pixel_data[56][48] = 0;
        pixel_data[56][49] = 0;
        pixel_data[56][50] = 0;
        pixel_data[56][51] = 0;
        pixel_data[56][52] = 0;
        pixel_data[56][53] = 0;
        pixel_data[56][54] = 0;
        pixel_data[56][55] = 0;
        pixel_data[56][56] = 0;
        pixel_data[56][57] = 0;
        pixel_data[56][58] = 0;
        pixel_data[56][59] = 0;
        pixel_data[56][60] = 0;
        pixel_data[56][61] = 0;
        pixel_data[56][62] = 0;
        pixel_data[56][63] = 0;
        pixel_data[56][64] = 0;
        pixel_data[56][65] = 0;
        pixel_data[56][66] = 0;
        pixel_data[56][67] = 0;
        pixel_data[56][68] = 0;
        pixel_data[56][69] = 0;
        pixel_data[56][70] = 0;
        pixel_data[56][71] = 0;
        pixel_data[56][72] = 0;
        pixel_data[56][73] = 0;
        pixel_data[56][74] = 0;
        pixel_data[56][75] = 0;
        pixel_data[56][76] = 0;
        pixel_data[56][77] = 0;
        pixel_data[56][78] = 0;
        pixel_data[56][79] = 0;
        pixel_data[56][80] = 0;
        pixel_data[56][81] = 0;
        pixel_data[56][82] = 0;
        pixel_data[56][83] = 0;
        pixel_data[56][84] = 0;
        pixel_data[56][85] = 0;
        pixel_data[56][86] = 0;
        pixel_data[56][87] = 0;
        pixel_data[56][88] = 0;
        pixel_data[56][89] = 0;
        pixel_data[56][90] = 0;
        pixel_data[56][91] = 0;
        pixel_data[56][92] = 0;
        pixel_data[56][93] = 0;
        pixel_data[56][94] = 0;
        pixel_data[56][95] = 0;
        pixel_data[56][96] = 0;
        pixel_data[56][97] = 0;
        pixel_data[56][98] = 0;
        pixel_data[56][99] = 0;
        pixel_data[56][100] = 0;
        pixel_data[56][101] = 0;
        pixel_data[56][102] = 0;
        pixel_data[56][103] = 0;
        pixel_data[56][104] = 0;
        pixel_data[56][105] = 0;
        pixel_data[56][106] = 0;
        pixel_data[56][107] = 0;
        pixel_data[56][108] = 0;
        pixel_data[56][109] = 0;
        pixel_data[56][110] = 0;
        pixel_data[56][111] = 0;
        pixel_data[56][112] = 0;
        pixel_data[56][113] = 0;
        pixel_data[56][114] = 0;
        pixel_data[56][115] = 0;
        pixel_data[56][116] = 0;
        pixel_data[56][117] = 0;
        pixel_data[56][118] = 0;
        pixel_data[56][119] = 0;
        pixel_data[56][120] = 0;
        pixel_data[56][121] = 0;
        pixel_data[56][122] = 0;
        pixel_data[56][123] = 0;
        pixel_data[56][124] = 0;
        pixel_data[56][125] = 0;
        pixel_data[56][126] = 0;
        pixel_data[56][127] = 0;
        pixel_data[56][128] = 0;
        pixel_data[56][129] = 0;
        pixel_data[56][130] = 0;
        pixel_data[56][131] = 0;
        pixel_data[56][132] = 0;
        pixel_data[56][133] = 0;
        pixel_data[56][134] = 0;
        pixel_data[56][135] = 0;
        pixel_data[56][136] = 0;
        pixel_data[56][137] = 0;
        pixel_data[56][138] = 0;
        pixel_data[56][139] = 0;
        pixel_data[56][140] = 0;
        pixel_data[56][141] = 0;
        pixel_data[56][142] = 0;
        pixel_data[56][143] = 0;
        pixel_data[56][144] = 0;
        pixel_data[56][145] = 0;
        pixel_data[56][146] = 0;
        pixel_data[56][147] = 0;
        pixel_data[56][148] = 0;
        pixel_data[56][149] = 0;
        pixel_data[56][150] = 0;
        pixel_data[56][151] = 0;
        pixel_data[56][152] = 0;
        pixel_data[56][153] = 0;
        pixel_data[56][154] = 0;
        pixel_data[56][155] = 0;
        pixel_data[56][156] = 0;
        pixel_data[56][157] = 0;
        pixel_data[56][158] = 0;
        pixel_data[56][159] = 0;
        pixel_data[56][160] = 0;
        pixel_data[56][161] = 0;
        pixel_data[56][162] = 0;
        pixel_data[56][163] = 0;
        pixel_data[56][164] = 0;
        pixel_data[56][165] = 0;
        pixel_data[56][166] = 0;
        pixel_data[56][167] = 0;
        pixel_data[56][168] = 0;
        pixel_data[56][169] = 0;
        pixel_data[56][170] = 0;
        pixel_data[56][171] = 0;
        pixel_data[56][172] = 0;
        pixel_data[56][173] = 0;
        pixel_data[56][174] = 0;
        pixel_data[56][175] = 0;
        pixel_data[56][176] = 0;
        pixel_data[56][177] = 0;
        pixel_data[56][178] = 0;
        pixel_data[56][179] = 0;
        pixel_data[56][180] = 0;
        pixel_data[56][181] = 0;
        pixel_data[56][182] = 0;
        pixel_data[56][183] = 0;
        pixel_data[56][184] = 0;
        pixel_data[56][185] = 0;
        pixel_data[56][186] = 0;
        pixel_data[56][187] = 0;
        pixel_data[56][188] = 0;
        pixel_data[56][189] = 0;
        pixel_data[56][190] = 0;
        pixel_data[56][191] = 0;
        pixel_data[56][192] = 0;
        pixel_data[56][193] = 0;
        pixel_data[56][194] = 0;
        pixel_data[56][195] = 0;
        pixel_data[56][196] = 0;
        pixel_data[56][197] = 0;
        pixel_data[56][198] = 0;
        pixel_data[56][199] = 0; // y=56
        pixel_data[57][0] = 0;
        pixel_data[57][1] = 0;
        pixel_data[57][2] = 0;
        pixel_data[57][3] = 0;
        pixel_data[57][4] = 0;
        pixel_data[57][5] = 0;
        pixel_data[57][6] = 0;
        pixel_data[57][7] = 0;
        pixel_data[57][8] = 0;
        pixel_data[57][9] = 0;
        pixel_data[57][10] = 0;
        pixel_data[57][11] = 0;
        pixel_data[57][12] = 0;
        pixel_data[57][13] = 0;
        pixel_data[57][14] = 0;
        pixel_data[57][15] = 0;
        pixel_data[57][16] = 0;
        pixel_data[57][17] = 0;
        pixel_data[57][18] = 0;
        pixel_data[57][19] = 0;
        pixel_data[57][20] = 0;
        pixel_data[57][21] = 0;
        pixel_data[57][22] = 0;
        pixel_data[57][23] = 0;
        pixel_data[57][24] = 0;
        pixel_data[57][25] = 0;
        pixel_data[57][26] = 0;
        pixel_data[57][27] = 0;
        pixel_data[57][28] = 0;
        pixel_data[57][29] = 0;
        pixel_data[57][30] = 0;
        pixel_data[57][31] = 0;
        pixel_data[57][32] = 0;
        pixel_data[57][33] = 0;
        pixel_data[57][34] = 0;
        pixel_data[57][35] = 0;
        pixel_data[57][36] = 0;
        pixel_data[57][37] = 0;
        pixel_data[57][38] = 0;
        pixel_data[57][39] = 0;
        pixel_data[57][40] = 0;
        pixel_data[57][41] = 0;
        pixel_data[57][42] = 0;
        pixel_data[57][43] = 0;
        pixel_data[57][44] = 0;
        pixel_data[57][45] = 0;
        pixel_data[57][46] = 0;
        pixel_data[57][47] = 0;
        pixel_data[57][48] = 0;
        pixel_data[57][49] = 0;
        pixel_data[57][50] = 0;
        pixel_data[57][51] = 0;
        pixel_data[57][52] = 0;
        pixel_data[57][53] = 0;
        pixel_data[57][54] = 0;
        pixel_data[57][55] = 0;
        pixel_data[57][56] = 0;
        pixel_data[57][57] = 0;
        pixel_data[57][58] = 0;
        pixel_data[57][59] = 0;
        pixel_data[57][60] = 0;
        pixel_data[57][61] = 0;
        pixel_data[57][62] = 0;
        pixel_data[57][63] = 0;
        pixel_data[57][64] = 0;
        pixel_data[57][65] = 0;
        pixel_data[57][66] = 0;
        pixel_data[57][67] = 0;
        pixel_data[57][68] = 0;
        pixel_data[57][69] = 0;
        pixel_data[57][70] = 0;
        pixel_data[57][71] = 0;
        pixel_data[57][72] = 0;
        pixel_data[57][73] = 0;
        pixel_data[57][74] = 0;
        pixel_data[57][75] = 0;
        pixel_data[57][76] = 0;
        pixel_data[57][77] = 0;
        pixel_data[57][78] = 0;
        pixel_data[57][79] = 0;
        pixel_data[57][80] = 0;
        pixel_data[57][81] = 0;
        pixel_data[57][82] = 0;
        pixel_data[57][83] = 0;
        pixel_data[57][84] = 0;
        pixel_data[57][85] = 0;
        pixel_data[57][86] = 0;
        pixel_data[57][87] = 0;
        pixel_data[57][88] = 0;
        pixel_data[57][89] = 0;
        pixel_data[57][90] = 0;
        pixel_data[57][91] = 0;
        pixel_data[57][92] = 0;
        pixel_data[57][93] = 0;
        pixel_data[57][94] = 0;
        pixel_data[57][95] = 0;
        pixel_data[57][96] = 0;
        pixel_data[57][97] = 0;
        pixel_data[57][98] = 0;
        pixel_data[57][99] = 0;
        pixel_data[57][100] = 0;
        pixel_data[57][101] = 0;
        pixel_data[57][102] = 0;
        pixel_data[57][103] = 0;
        pixel_data[57][104] = 0;
        pixel_data[57][105] = 0;
        pixel_data[57][106] = 0;
        pixel_data[57][107] = 0;
        pixel_data[57][108] = 0;
        pixel_data[57][109] = 0;
        pixel_data[57][110] = 0;
        pixel_data[57][111] = 0;
        pixel_data[57][112] = 0;
        pixel_data[57][113] = 0;
        pixel_data[57][114] = 0;
        pixel_data[57][115] = 0;
        pixel_data[57][116] = 0;
        pixel_data[57][117] = 0;
        pixel_data[57][118] = 0;
        pixel_data[57][119] = 0;
        pixel_data[57][120] = 0;
        pixel_data[57][121] = 0;
        pixel_data[57][122] = 0;
        pixel_data[57][123] = 0;
        pixel_data[57][124] = 0;
        pixel_data[57][125] = 0;
        pixel_data[57][126] = 0;
        pixel_data[57][127] = 0;
        pixel_data[57][128] = 0;
        pixel_data[57][129] = 0;
        pixel_data[57][130] = 0;
        pixel_data[57][131] = 0;
        pixel_data[57][132] = 0;
        pixel_data[57][133] = 0;
        pixel_data[57][134] = 0;
        pixel_data[57][135] = 0;
        pixel_data[57][136] = 0;
        pixel_data[57][137] = 0;
        pixel_data[57][138] = 0;
        pixel_data[57][139] = 0;
        pixel_data[57][140] = 0;
        pixel_data[57][141] = 0;
        pixel_data[57][142] = 0;
        pixel_data[57][143] = 0;
        pixel_data[57][144] = 0;
        pixel_data[57][145] = 0;
        pixel_data[57][146] = 0;
        pixel_data[57][147] = 0;
        pixel_data[57][148] = 0;
        pixel_data[57][149] = 0;
        pixel_data[57][150] = 0;
        pixel_data[57][151] = 0;
        pixel_data[57][152] = 0;
        pixel_data[57][153] = 0;
        pixel_data[57][154] = 0;
        pixel_data[57][155] = 0;
        pixel_data[57][156] = 0;
        pixel_data[57][157] = 0;
        pixel_data[57][158] = 0;
        pixel_data[57][159] = 0;
        pixel_data[57][160] = 0;
        pixel_data[57][161] = 0;
        pixel_data[57][162] = 0;
        pixel_data[57][163] = 0;
        pixel_data[57][164] = 0;
        pixel_data[57][165] = 0;
        pixel_data[57][166] = 0;
        pixel_data[57][167] = 0;
        pixel_data[57][168] = 0;
        pixel_data[57][169] = 0;
        pixel_data[57][170] = 0;
        pixel_data[57][171] = 0;
        pixel_data[57][172] = 0;
        pixel_data[57][173] = 0;
        pixel_data[57][174] = 0;
        pixel_data[57][175] = 0;
        pixel_data[57][176] = 0;
        pixel_data[57][177] = 0;
        pixel_data[57][178] = 0;
        pixel_data[57][179] = 0;
        pixel_data[57][180] = 0;
        pixel_data[57][181] = 0;
        pixel_data[57][182] = 0;
        pixel_data[57][183] = 0;
        pixel_data[57][184] = 0;
        pixel_data[57][185] = 0;
        pixel_data[57][186] = 0;
        pixel_data[57][187] = 0;
        pixel_data[57][188] = 0;
        pixel_data[57][189] = 0;
        pixel_data[57][190] = 0;
        pixel_data[57][191] = 0;
        pixel_data[57][192] = 0;
        pixel_data[57][193] = 0;
        pixel_data[57][194] = 0;
        pixel_data[57][195] = 0;
        pixel_data[57][196] = 0;
        pixel_data[57][197] = 0;
        pixel_data[57][198] = 0;
        pixel_data[57][199] = 0; // y=57
        pixel_data[58][0] = 0;
        pixel_data[58][1] = 0;
        pixel_data[58][2] = 0;
        pixel_data[58][3] = 0;
        pixel_data[58][4] = 0;
        pixel_data[58][5] = 0;
        pixel_data[58][6] = 0;
        pixel_data[58][7] = 0;
        pixel_data[58][8] = 0;
        pixel_data[58][9] = 0;
        pixel_data[58][10] = 0;
        pixel_data[58][11] = 0;
        pixel_data[58][12] = 0;
        pixel_data[58][13] = 0;
        pixel_data[58][14] = 0;
        pixel_data[58][15] = 0;
        pixel_data[58][16] = 0;
        pixel_data[58][17] = 0;
        pixel_data[58][18] = 0;
        pixel_data[58][19] = 0;
        pixel_data[58][20] = 0;
        pixel_data[58][21] = 0;
        pixel_data[58][22] = 0;
        pixel_data[58][23] = 0;
        pixel_data[58][24] = 0;
        pixel_data[58][25] = 0;
        pixel_data[58][26] = 0;
        pixel_data[58][27] = 0;
        pixel_data[58][28] = 0;
        pixel_data[58][29] = 0;
        pixel_data[58][30] = 0;
        pixel_data[58][31] = 0;
        pixel_data[58][32] = 0;
        pixel_data[58][33] = 0;
        pixel_data[58][34] = 0;
        pixel_data[58][35] = 0;
        pixel_data[58][36] = 0;
        pixel_data[58][37] = 0;
        pixel_data[58][38] = 0;
        pixel_data[58][39] = 0;
        pixel_data[58][40] = 0;
        pixel_data[58][41] = 0;
        pixel_data[58][42] = 0;
        pixel_data[58][43] = 0;
        pixel_data[58][44] = 0;
        pixel_data[58][45] = 0;
        pixel_data[58][46] = 0;
        pixel_data[58][47] = 0;
        pixel_data[58][48] = 0;
        pixel_data[58][49] = 0;
        pixel_data[58][50] = 0;
        pixel_data[58][51] = 0;
        pixel_data[58][52] = 0;
        pixel_data[58][53] = 0;
        pixel_data[58][54] = 0;
        pixel_data[58][55] = 0;
        pixel_data[58][56] = 0;
        pixel_data[58][57] = 0;
        pixel_data[58][58] = 0;
        pixel_data[58][59] = 0;
        pixel_data[58][60] = 0;
        pixel_data[58][61] = 0;
        pixel_data[58][62] = 0;
        pixel_data[58][63] = 0;
        pixel_data[58][64] = 0;
        pixel_data[58][65] = 0;
        pixel_data[58][66] = 0;
        pixel_data[58][67] = 0;
        pixel_data[58][68] = 0;
        pixel_data[58][69] = 0;
        pixel_data[58][70] = 0;
        pixel_data[58][71] = 0;
        pixel_data[58][72] = 0;
        pixel_data[58][73] = 0;
        pixel_data[58][74] = 0;
        pixel_data[58][75] = 0;
        pixel_data[58][76] = 0;
        pixel_data[58][77] = 0;
        pixel_data[58][78] = 0;
        pixel_data[58][79] = 0;
        pixel_data[58][80] = 0;
        pixel_data[58][81] = 0;
        pixel_data[58][82] = 0;
        pixel_data[58][83] = 0;
        pixel_data[58][84] = 0;
        pixel_data[58][85] = 0;
        pixel_data[58][86] = 0;
        pixel_data[58][87] = 0;
        pixel_data[58][88] = 0;
        pixel_data[58][89] = 0;
        pixel_data[58][90] = 0;
        pixel_data[58][91] = 0;
        pixel_data[58][92] = 0;
        pixel_data[58][93] = 0;
        pixel_data[58][94] = 0;
        pixel_data[58][95] = 0;
        pixel_data[58][96] = 0;
        pixel_data[58][97] = 0;
        pixel_data[58][98] = 0;
        pixel_data[58][99] = 0;
        pixel_data[58][100] = 0;
        pixel_data[58][101] = 0;
        pixel_data[58][102] = 0;
        pixel_data[58][103] = 0;
        pixel_data[58][104] = 0;
        pixel_data[58][105] = 0;
        pixel_data[58][106] = 0;
        pixel_data[58][107] = 0;
        pixel_data[58][108] = 0;
        pixel_data[58][109] = 0;
        pixel_data[58][110] = 0;
        pixel_data[58][111] = 0;
        pixel_data[58][112] = 0;
        pixel_data[58][113] = 0;
        pixel_data[58][114] = 0;
        pixel_data[58][115] = 0;
        pixel_data[58][116] = 0;
        pixel_data[58][117] = 0;
        pixel_data[58][118] = 0;
        pixel_data[58][119] = 0;
        pixel_data[58][120] = 0;
        pixel_data[58][121] = 0;
        pixel_data[58][122] = 0;
        pixel_data[58][123] = 0;
        pixel_data[58][124] = 0;
        pixel_data[58][125] = 0;
        pixel_data[58][126] = 0;
        pixel_data[58][127] = 0;
        pixel_data[58][128] = 0;
        pixel_data[58][129] = 0;
        pixel_data[58][130] = 0;
        pixel_data[58][131] = 0;
        pixel_data[58][132] = 0;
        pixel_data[58][133] = 0;
        pixel_data[58][134] = 0;
        pixel_data[58][135] = 0;
        pixel_data[58][136] = 0;
        pixel_data[58][137] = 0;
        pixel_data[58][138] = 0;
        pixel_data[58][139] = 0;
        pixel_data[58][140] = 0;
        pixel_data[58][141] = 0;
        pixel_data[58][142] = 0;
        pixel_data[58][143] = 0;
        pixel_data[58][144] = 0;
        pixel_data[58][145] = 0;
        pixel_data[58][146] = 0;
        pixel_data[58][147] = 0;
        pixel_data[58][148] = 0;
        pixel_data[58][149] = 0;
        pixel_data[58][150] = 0;
        pixel_data[58][151] = 0;
        pixel_data[58][152] = 0;
        pixel_data[58][153] = 0;
        pixel_data[58][154] = 0;
        pixel_data[58][155] = 0;
        pixel_data[58][156] = 0;
        pixel_data[58][157] = 0;
        pixel_data[58][158] = 0;
        pixel_data[58][159] = 0;
        pixel_data[58][160] = 0;
        pixel_data[58][161] = 0;
        pixel_data[58][162] = 0;
        pixel_data[58][163] = 0;
        pixel_data[58][164] = 0;
        pixel_data[58][165] = 0;
        pixel_data[58][166] = 0;
        pixel_data[58][167] = 0;
        pixel_data[58][168] = 0;
        pixel_data[58][169] = 0;
        pixel_data[58][170] = 0;
        pixel_data[58][171] = 0;
        pixel_data[58][172] = 0;
        pixel_data[58][173] = 0;
        pixel_data[58][174] = 0;
        pixel_data[58][175] = 0;
        pixel_data[58][176] = 0;
        pixel_data[58][177] = 0;
        pixel_data[58][178] = 0;
        pixel_data[58][179] = 0;
        pixel_data[58][180] = 0;
        pixel_data[58][181] = 0;
        pixel_data[58][182] = 0;
        pixel_data[58][183] = 0;
        pixel_data[58][184] = 0;
        pixel_data[58][185] = 0;
        pixel_data[58][186] = 0;
        pixel_data[58][187] = 0;
        pixel_data[58][188] = 0;
        pixel_data[58][189] = 0;
        pixel_data[58][190] = 0;
        pixel_data[58][191] = 0;
        pixel_data[58][192] = 0;
        pixel_data[58][193] = 0;
        pixel_data[58][194] = 0;
        pixel_data[58][195] = 0;
        pixel_data[58][196] = 0;
        pixel_data[58][197] = 0;
        pixel_data[58][198] = 0;
        pixel_data[58][199] = 0; // y=58
        pixel_data[59][0] = 0;
        pixel_data[59][1] = 0;
        pixel_data[59][2] = 0;
        pixel_data[59][3] = 0;
        pixel_data[59][4] = 0;
        pixel_data[59][5] = 0;
        pixel_data[59][6] = 0;
        pixel_data[59][7] = 0;
        pixel_data[59][8] = 0;
        pixel_data[59][9] = 0;
        pixel_data[59][10] = 0;
        pixel_data[59][11] = 0;
        pixel_data[59][12] = 0;
        pixel_data[59][13] = 0;
        pixel_data[59][14] = 0;
        pixel_data[59][15] = 0;
        pixel_data[59][16] = 0;
        pixel_data[59][17] = 0;
        pixel_data[59][18] = 0;
        pixel_data[59][19] = 0;
        pixel_data[59][20] = 0;
        pixel_data[59][21] = 0;
        pixel_data[59][22] = 0;
        pixel_data[59][23] = 0;
        pixel_data[59][24] = 0;
        pixel_data[59][25] = 0;
        pixel_data[59][26] = 0;
        pixel_data[59][27] = 0;
        pixel_data[59][28] = 0;
        pixel_data[59][29] = 0;
        pixel_data[59][30] = 0;
        pixel_data[59][31] = 0;
        pixel_data[59][32] = 0;
        pixel_data[59][33] = 0;
        pixel_data[59][34] = 0;
        pixel_data[59][35] = 0;
        pixel_data[59][36] = 0;
        pixel_data[59][37] = 0;
        pixel_data[59][38] = 0;
        pixel_data[59][39] = 0;
        pixel_data[59][40] = 0;
        pixel_data[59][41] = 0;
        pixel_data[59][42] = 0;
        pixel_data[59][43] = 0;
        pixel_data[59][44] = 0;
        pixel_data[59][45] = 0;
        pixel_data[59][46] = 0;
        pixel_data[59][47] = 0;
        pixel_data[59][48] = 0;
        pixel_data[59][49] = 0;
        pixel_data[59][50] = 0;
        pixel_data[59][51] = 0;
        pixel_data[59][52] = 0;
        pixel_data[59][53] = 0;
        pixel_data[59][54] = 0;
        pixel_data[59][55] = 0;
        pixel_data[59][56] = 0;
        pixel_data[59][57] = 0;
        pixel_data[59][58] = 0;
        pixel_data[59][59] = 0;
        pixel_data[59][60] = 0;
        pixel_data[59][61] = 0;
        pixel_data[59][62] = 0;
        pixel_data[59][63] = 0;
        pixel_data[59][64] = 0;
        pixel_data[59][65] = 0;
        pixel_data[59][66] = 0;
        pixel_data[59][67] = 0;
        pixel_data[59][68] = 0;
        pixel_data[59][69] = 0;
        pixel_data[59][70] = 0;
        pixel_data[59][71] = 0;
        pixel_data[59][72] = 0;
        pixel_data[59][73] = 0;
        pixel_data[59][74] = 0;
        pixel_data[59][75] = 0;
        pixel_data[59][76] = 0;
        pixel_data[59][77] = 0;
        pixel_data[59][78] = 0;
        pixel_data[59][79] = 0;
        pixel_data[59][80] = 0;
        pixel_data[59][81] = 0;
        pixel_data[59][82] = 0;
        pixel_data[59][83] = 0;
        pixel_data[59][84] = 0;
        pixel_data[59][85] = 0;
        pixel_data[59][86] = 0;
        pixel_data[59][87] = 0;
        pixel_data[59][88] = 0;
        pixel_data[59][89] = 0;
        pixel_data[59][90] = 0;
        pixel_data[59][91] = 0;
        pixel_data[59][92] = 0;
        pixel_data[59][93] = 0;
        pixel_data[59][94] = 0;
        pixel_data[59][95] = 0;
        pixel_data[59][96] = 0;
        pixel_data[59][97] = 0;
        pixel_data[59][98] = 0;
        pixel_data[59][99] = 0;
        pixel_data[59][100] = 0;
        pixel_data[59][101] = 0;
        pixel_data[59][102] = 0;
        pixel_data[59][103] = 0;
        pixel_data[59][104] = 0;
        pixel_data[59][105] = 0;
        pixel_data[59][106] = 0;
        pixel_data[59][107] = 0;
        pixel_data[59][108] = 0;
        pixel_data[59][109] = 0;
        pixel_data[59][110] = 0;
        pixel_data[59][111] = 0;
        pixel_data[59][112] = 0;
        pixel_data[59][113] = 0;
        pixel_data[59][114] = 0;
        pixel_data[59][115] = 0;
        pixel_data[59][116] = 0;
        pixel_data[59][117] = 0;
        pixel_data[59][118] = 0;
        pixel_data[59][119] = 0;
        pixel_data[59][120] = 0;
        pixel_data[59][121] = 0;
        pixel_data[59][122] = 0;
        pixel_data[59][123] = 0;
        pixel_data[59][124] = 0;
        pixel_data[59][125] = 0;
        pixel_data[59][126] = 0;
        pixel_data[59][127] = 0;
        pixel_data[59][128] = 0;
        pixel_data[59][129] = 0;
        pixel_data[59][130] = 0;
        pixel_data[59][131] = 0;
        pixel_data[59][132] = 0;
        pixel_data[59][133] = 0;
        pixel_data[59][134] = 0;
        pixel_data[59][135] = 0;
        pixel_data[59][136] = 0;
        pixel_data[59][137] = 0;
        pixel_data[59][138] = 0;
        pixel_data[59][139] = 0;
        pixel_data[59][140] = 0;
        pixel_data[59][141] = 0;
        pixel_data[59][142] = 0;
        pixel_data[59][143] = 0;
        pixel_data[59][144] = 0;
        pixel_data[59][145] = 0;
        pixel_data[59][146] = 0;
        pixel_data[59][147] = 0;
        pixel_data[59][148] = 0;
        pixel_data[59][149] = 0;
        pixel_data[59][150] = 0;
        pixel_data[59][151] = 0;
        pixel_data[59][152] = 0;
        pixel_data[59][153] = 0;
        pixel_data[59][154] = 0;
        pixel_data[59][155] = 0;
        pixel_data[59][156] = 0;
        pixel_data[59][157] = 0;
        pixel_data[59][158] = 0;
        pixel_data[59][159] = 0;
        pixel_data[59][160] = 0;
        pixel_data[59][161] = 0;
        pixel_data[59][162] = 0;
        pixel_data[59][163] = 0;
        pixel_data[59][164] = 0;
        pixel_data[59][165] = 0;
        pixel_data[59][166] = 0;
        pixel_data[59][167] = 0;
        pixel_data[59][168] = 0;
        pixel_data[59][169] = 0;
        pixel_data[59][170] = 0;
        pixel_data[59][171] = 0;
        pixel_data[59][172] = 0;
        pixel_data[59][173] = 0;
        pixel_data[59][174] = 0;
        pixel_data[59][175] = 0;
        pixel_data[59][176] = 0;
        pixel_data[59][177] = 0;
        pixel_data[59][178] = 0;
        pixel_data[59][179] = 0;
        pixel_data[59][180] = 0;
        pixel_data[59][181] = 0;
        pixel_data[59][182] = 0;
        pixel_data[59][183] = 0;
        pixel_data[59][184] = 0;
        pixel_data[59][185] = 0;
        pixel_data[59][186] = 0;
        pixel_data[59][187] = 0;
        pixel_data[59][188] = 0;
        pixel_data[59][189] = 0;
        pixel_data[59][190] = 0;
        pixel_data[59][191] = 0;
        pixel_data[59][192] = 0;
        pixel_data[59][193] = 0;
        pixel_data[59][194] = 0;
        pixel_data[59][195] = 0;
        pixel_data[59][196] = 0;
        pixel_data[59][197] = 0;
        pixel_data[59][198] = 0;
        pixel_data[59][199] = 0; // y=59
        pixel_data[60][0] = 0;
        pixel_data[60][1] = 0;
        pixel_data[60][2] = 0;
        pixel_data[60][3] = 0;
        pixel_data[60][4] = 0;
        pixel_data[60][5] = 0;
        pixel_data[60][6] = 0;
        pixel_data[60][7] = 0;
        pixel_data[60][8] = 0;
        pixel_data[60][9] = 0;
        pixel_data[60][10] = 0;
        pixel_data[60][11] = 0;
        pixel_data[60][12] = 0;
        pixel_data[60][13] = 0;
        pixel_data[60][14] = 0;
        pixel_data[60][15] = 0;
        pixel_data[60][16] = 0;
        pixel_data[60][17] = 0;
        pixel_data[60][18] = 0;
        pixel_data[60][19] = 0;
        pixel_data[60][20] = 0;
        pixel_data[60][21] = 0;
        pixel_data[60][22] = 0;
        pixel_data[60][23] = 0;
        pixel_data[60][24] = 0;
        pixel_data[60][25] = 0;
        pixel_data[60][26] = 0;
        pixel_data[60][27] = 0;
        pixel_data[60][28] = 0;
        pixel_data[60][29] = 0;
        pixel_data[60][30] = 0;
        pixel_data[60][31] = 0;
        pixel_data[60][32] = 0;
        pixel_data[60][33] = 0;
        pixel_data[60][34] = 0;
        pixel_data[60][35] = 0;
        pixel_data[60][36] = 0;
        pixel_data[60][37] = 0;
        pixel_data[60][38] = 0;
        pixel_data[60][39] = 0;
        pixel_data[60][40] = 0;
        pixel_data[60][41] = 0;
        pixel_data[60][42] = 0;
        pixel_data[60][43] = 0;
        pixel_data[60][44] = 0;
        pixel_data[60][45] = 0;
        pixel_data[60][46] = 0;
        pixel_data[60][47] = 0;
        pixel_data[60][48] = 0;
        pixel_data[60][49] = 0;
        pixel_data[60][50] = 0;
        pixel_data[60][51] = 0;
        pixel_data[60][52] = 0;
        pixel_data[60][53] = 0;
        pixel_data[60][54] = 0;
        pixel_data[60][55] = 0;
        pixel_data[60][56] = 0;
        pixel_data[60][57] = 0;
        pixel_data[60][58] = 0;
        pixel_data[60][59] = 0;
        pixel_data[60][60] = 0;
        pixel_data[60][61] = 0;
        pixel_data[60][62] = 0;
        pixel_data[60][63] = 0;
        pixel_data[60][64] = 0;
        pixel_data[60][65] = 0;
        pixel_data[60][66] = 0;
        pixel_data[60][67] = 0;
        pixel_data[60][68] = 0;
        pixel_data[60][69] = 0;
        pixel_data[60][70] = 0;
        pixel_data[60][71] = 0;
        pixel_data[60][72] = 0;
        pixel_data[60][73] = 0;
        pixel_data[60][74] = 0;
        pixel_data[60][75] = 0;
        pixel_data[60][76] = 0;
        pixel_data[60][77] = 0;
        pixel_data[60][78] = 0;
        pixel_data[60][79] = 0;
        pixel_data[60][80] = 0;
        pixel_data[60][81] = 0;
        pixel_data[60][82] = 0;
        pixel_data[60][83] = 0;
        pixel_data[60][84] = 0;
        pixel_data[60][85] = 0;
        pixel_data[60][86] = 0;
        pixel_data[60][87] = 0;
        pixel_data[60][88] = 0;
        pixel_data[60][89] = 0;
        pixel_data[60][90] = 0;
        pixel_data[60][91] = 0;
        pixel_data[60][92] = 0;
        pixel_data[60][93] = 0;
        pixel_data[60][94] = 0;
        pixel_data[60][95] = 0;
        pixel_data[60][96] = 0;
        pixel_data[60][97] = 0;
        pixel_data[60][98] = 0;
        pixel_data[60][99] = 0;
        pixel_data[60][100] = 0;
        pixel_data[60][101] = 0;
        pixel_data[60][102] = 0;
        pixel_data[60][103] = 0;
        pixel_data[60][104] = 0;
        pixel_data[60][105] = 0;
        pixel_data[60][106] = 0;
        pixel_data[60][107] = 0;
        pixel_data[60][108] = 0;
        pixel_data[60][109] = 0;
        pixel_data[60][110] = 0;
        pixel_data[60][111] = 0;
        pixel_data[60][112] = 0;
        pixel_data[60][113] = 0;
        pixel_data[60][114] = 0;
        pixel_data[60][115] = 0;
        pixel_data[60][116] = 0;
        pixel_data[60][117] = 0;
        pixel_data[60][118] = 0;
        pixel_data[60][119] = 0;
        pixel_data[60][120] = 0;
        pixel_data[60][121] = 0;
        pixel_data[60][122] = 0;
        pixel_data[60][123] = 0;
        pixel_data[60][124] = 0;
        pixel_data[60][125] = 0;
        pixel_data[60][126] = 0;
        pixel_data[60][127] = 0;
        pixel_data[60][128] = 0;
        pixel_data[60][129] = 0;
        pixel_data[60][130] = 0;
        pixel_data[60][131] = 0;
        pixel_data[60][132] = 0;
        pixel_data[60][133] = 0;
        pixel_data[60][134] = 0;
        pixel_data[60][135] = 0;
        pixel_data[60][136] = 0;
        pixel_data[60][137] = 0;
        pixel_data[60][138] = 0;
        pixel_data[60][139] = 0;
        pixel_data[60][140] = 0;
        pixel_data[60][141] = 0;
        pixel_data[60][142] = 0;
        pixel_data[60][143] = 0;
        pixel_data[60][144] = 0;
        pixel_data[60][145] = 0;
        pixel_data[60][146] = 0;
        pixel_data[60][147] = 0;
        pixel_data[60][148] = 0;
        pixel_data[60][149] = 0;
        pixel_data[60][150] = 0;
        pixel_data[60][151] = 0;
        pixel_data[60][152] = 0;
        pixel_data[60][153] = 0;
        pixel_data[60][154] = 0;
        pixel_data[60][155] = 0;
        pixel_data[60][156] = 0;
        pixel_data[60][157] = 0;
        pixel_data[60][158] = 0;
        pixel_data[60][159] = 0;
        pixel_data[60][160] = 0;
        pixel_data[60][161] = 0;
        pixel_data[60][162] = 0;
        pixel_data[60][163] = 0;
        pixel_data[60][164] = 0;
        pixel_data[60][165] = 0;
        pixel_data[60][166] = 0;
        pixel_data[60][167] = 0;
        pixel_data[60][168] = 0;
        pixel_data[60][169] = 0;
        pixel_data[60][170] = 0;
        pixel_data[60][171] = 0;
        pixel_data[60][172] = 0;
        pixel_data[60][173] = 0;
        pixel_data[60][174] = 0;
        pixel_data[60][175] = 0;
        pixel_data[60][176] = 0;
        pixel_data[60][177] = 0;
        pixel_data[60][178] = 0;
        pixel_data[60][179] = 0;
        pixel_data[60][180] = 0;
        pixel_data[60][181] = 0;
        pixel_data[60][182] = 0;
        pixel_data[60][183] = 0;
        pixel_data[60][184] = 0;
        pixel_data[60][185] = 0;
        pixel_data[60][186] = 0;
        pixel_data[60][187] = 0;
        pixel_data[60][188] = 0;
        pixel_data[60][189] = 0;
        pixel_data[60][190] = 0;
        pixel_data[60][191] = 0;
        pixel_data[60][192] = 0;
        pixel_data[60][193] = 0;
        pixel_data[60][194] = 0;
        pixel_data[60][195] = 0;
        pixel_data[60][196] = 0;
        pixel_data[60][197] = 0;
        pixel_data[60][198] = 0;
        pixel_data[60][199] = 0; // y=60
        pixel_data[61][0] = 0;
        pixel_data[61][1] = 0;
        pixel_data[61][2] = 0;
        pixel_data[61][3] = 0;
        pixel_data[61][4] = 0;
        pixel_data[61][5] = 0;
        pixel_data[61][6] = 0;
        pixel_data[61][7] = 0;
        pixel_data[61][8] = 0;
        pixel_data[61][9] = 0;
        pixel_data[61][10] = 0;
        pixel_data[61][11] = 0;
        pixel_data[61][12] = 0;
        pixel_data[61][13] = 0;
        pixel_data[61][14] = 0;
        pixel_data[61][15] = 0;
        pixel_data[61][16] = 0;
        pixel_data[61][17] = 0;
        pixel_data[61][18] = 0;
        pixel_data[61][19] = 0;
        pixel_data[61][20] = 0;
        pixel_data[61][21] = 0;
        pixel_data[61][22] = 0;
        pixel_data[61][23] = 0;
        pixel_data[61][24] = 0;
        pixel_data[61][25] = 0;
        pixel_data[61][26] = 0;
        pixel_data[61][27] = 0;
        pixel_data[61][28] = 0;
        pixel_data[61][29] = 0;
        pixel_data[61][30] = 0;
        pixel_data[61][31] = 0;
        pixel_data[61][32] = 0;
        pixel_data[61][33] = 0;
        pixel_data[61][34] = 0;
        pixel_data[61][35] = 0;
        pixel_data[61][36] = 0;
        pixel_data[61][37] = 0;
        pixel_data[61][38] = 0;
        pixel_data[61][39] = 0;
        pixel_data[61][40] = 0;
        pixel_data[61][41] = 0;
        pixel_data[61][42] = 0;
        pixel_data[61][43] = 0;
        pixel_data[61][44] = 0;
        pixel_data[61][45] = 0;
        pixel_data[61][46] = 0;
        pixel_data[61][47] = 0;
        pixel_data[61][48] = 0;
        pixel_data[61][49] = 0;
        pixel_data[61][50] = 0;
        pixel_data[61][51] = 0;
        pixel_data[61][52] = 0;
        pixel_data[61][53] = 0;
        pixel_data[61][54] = 0;
        pixel_data[61][55] = 0;
        pixel_data[61][56] = 0;
        pixel_data[61][57] = 0;
        pixel_data[61][58] = 0;
        pixel_data[61][59] = 0;
        pixel_data[61][60] = 0;
        pixel_data[61][61] = 0;
        pixel_data[61][62] = 0;
        pixel_data[61][63] = 0;
        pixel_data[61][64] = 0;
        pixel_data[61][65] = 0;
        pixel_data[61][66] = 0;
        pixel_data[61][67] = 0;
        pixel_data[61][68] = 0;
        pixel_data[61][69] = 0;
        pixel_data[61][70] = 0;
        pixel_data[61][71] = 0;
        pixel_data[61][72] = 0;
        pixel_data[61][73] = 0;
        pixel_data[61][74] = 0;
        pixel_data[61][75] = 0;
        pixel_data[61][76] = 0;
        pixel_data[61][77] = 0;
        pixel_data[61][78] = 0;
        pixel_data[61][79] = 0;
        pixel_data[61][80] = 0;
        pixel_data[61][81] = 0;
        pixel_data[61][82] = 0;
        pixel_data[61][83] = 0;
        pixel_data[61][84] = 0;
        pixel_data[61][85] = 0;
        pixel_data[61][86] = 0;
        pixel_data[61][87] = 0;
        pixel_data[61][88] = 0;
        pixel_data[61][89] = 0;
        pixel_data[61][90] = 0;
        pixel_data[61][91] = 0;
        pixel_data[61][92] = 0;
        pixel_data[61][93] = 0;
        pixel_data[61][94] = 0;
        pixel_data[61][95] = 0;
        pixel_data[61][96] = 0;
        pixel_data[61][97] = 0;
        pixel_data[61][98] = 0;
        pixel_data[61][99] = 0;
        pixel_data[61][100] = 0;
        pixel_data[61][101] = 0;
        pixel_data[61][102] = 0;
        pixel_data[61][103] = 0;
        pixel_data[61][104] = 0;
        pixel_data[61][105] = 0;
        pixel_data[61][106] = 0;
        pixel_data[61][107] = 0;
        pixel_data[61][108] = 0;
        pixel_data[61][109] = 0;
        pixel_data[61][110] = 0;
        pixel_data[61][111] = 0;
        pixel_data[61][112] = 0;
        pixel_data[61][113] = 0;
        pixel_data[61][114] = 0;
        pixel_data[61][115] = 0;
        pixel_data[61][116] = 0;
        pixel_data[61][117] = 0;
        pixel_data[61][118] = 0;
        pixel_data[61][119] = 0;
        pixel_data[61][120] = 0;
        pixel_data[61][121] = 0;
        pixel_data[61][122] = 0;
        pixel_data[61][123] = 0;
        pixel_data[61][124] = 0;
        pixel_data[61][125] = 0;
        pixel_data[61][126] = 0;
        pixel_data[61][127] = 0;
        pixel_data[61][128] = 0;
        pixel_data[61][129] = 0;
        pixel_data[61][130] = 0;
        pixel_data[61][131] = 0;
        pixel_data[61][132] = 0;
        pixel_data[61][133] = 0;
        pixel_data[61][134] = 0;
        pixel_data[61][135] = 0;
        pixel_data[61][136] = 0;
        pixel_data[61][137] = 0;
        pixel_data[61][138] = 0;
        pixel_data[61][139] = 0;
        pixel_data[61][140] = 0;
        pixel_data[61][141] = 0;
        pixel_data[61][142] = 0;
        pixel_data[61][143] = 0;
        pixel_data[61][144] = 0;
        pixel_data[61][145] = 0;
        pixel_data[61][146] = 0;
        pixel_data[61][147] = 0;
        pixel_data[61][148] = 0;
        pixel_data[61][149] = 0;
        pixel_data[61][150] = 0;
        pixel_data[61][151] = 0;
        pixel_data[61][152] = 0;
        pixel_data[61][153] = 0;
        pixel_data[61][154] = 0;
        pixel_data[61][155] = 0;
        pixel_data[61][156] = 0;
        pixel_data[61][157] = 0;
        pixel_data[61][158] = 0;
        pixel_data[61][159] = 0;
        pixel_data[61][160] = 0;
        pixel_data[61][161] = 0;
        pixel_data[61][162] = 0;
        pixel_data[61][163] = 0;
        pixel_data[61][164] = 0;
        pixel_data[61][165] = 0;
        pixel_data[61][166] = 0;
        pixel_data[61][167] = 0;
        pixel_data[61][168] = 0;
        pixel_data[61][169] = 0;
        pixel_data[61][170] = 0;
        pixel_data[61][171] = 0;
        pixel_data[61][172] = 0;
        pixel_data[61][173] = 0;
        pixel_data[61][174] = 0;
        pixel_data[61][175] = 0;
        pixel_data[61][176] = 0;
        pixel_data[61][177] = 0;
        pixel_data[61][178] = 0;
        pixel_data[61][179] = 0;
        pixel_data[61][180] = 0;
        pixel_data[61][181] = 0;
        pixel_data[61][182] = 0;
        pixel_data[61][183] = 0;
        pixel_data[61][184] = 0;
        pixel_data[61][185] = 0;
        pixel_data[61][186] = 0;
        pixel_data[61][187] = 0;
        pixel_data[61][188] = 0;
        pixel_data[61][189] = 0;
        pixel_data[61][190] = 0;
        pixel_data[61][191] = 0;
        pixel_data[61][192] = 0;
        pixel_data[61][193] = 0;
        pixel_data[61][194] = 0;
        pixel_data[61][195] = 0;
        pixel_data[61][196] = 0;
        pixel_data[61][197] = 0;
        pixel_data[61][198] = 0;
        pixel_data[61][199] = 0; // y=61
        pixel_data[62][0] = 0;
        pixel_data[62][1] = 0;
        pixel_data[62][2] = 0;
        pixel_data[62][3] = 0;
        pixel_data[62][4] = 0;
        pixel_data[62][5] = 0;
        pixel_data[62][6] = 0;
        pixel_data[62][7] = 0;
        pixel_data[62][8] = 0;
        pixel_data[62][9] = 0;
        pixel_data[62][10] = 0;
        pixel_data[62][11] = 0;
        pixel_data[62][12] = 0;
        pixel_data[62][13] = 0;
        pixel_data[62][14] = 0;
        pixel_data[62][15] = 0;
        pixel_data[62][16] = 0;
        pixel_data[62][17] = 0;
        pixel_data[62][18] = 0;
        pixel_data[62][19] = 0;
        pixel_data[62][20] = 0;
        pixel_data[62][21] = 0;
        pixel_data[62][22] = 0;
        pixel_data[62][23] = 0;
        pixel_data[62][24] = 0;
        pixel_data[62][25] = 0;
        pixel_data[62][26] = 0;
        pixel_data[62][27] = 0;
        pixel_data[62][28] = 0;
        pixel_data[62][29] = 0;
        pixel_data[62][30] = 0;
        pixel_data[62][31] = 0;
        pixel_data[62][32] = 0;
        pixel_data[62][33] = 0;
        pixel_data[62][34] = 0;
        pixel_data[62][35] = 0;
        pixel_data[62][36] = 0;
        pixel_data[62][37] = 0;
        pixel_data[62][38] = 0;
        pixel_data[62][39] = 0;
        pixel_data[62][40] = 0;
        pixel_data[62][41] = 0;
        pixel_data[62][42] = 0;
        pixel_data[62][43] = 0;
        pixel_data[62][44] = 0;
        pixel_data[62][45] = 0;
        pixel_data[62][46] = 0;
        pixel_data[62][47] = 0;
        pixel_data[62][48] = 0;
        pixel_data[62][49] = 0;
        pixel_data[62][50] = 0;
        pixel_data[62][51] = 0;
        pixel_data[62][52] = 0;
        pixel_data[62][53] = 0;
        pixel_data[62][54] = 0;
        pixel_data[62][55] = 0;
        pixel_data[62][56] = 0;
        pixel_data[62][57] = 0;
        pixel_data[62][58] = 0;
        pixel_data[62][59] = 0;
        pixel_data[62][60] = 0;
        pixel_data[62][61] = 0;
        pixel_data[62][62] = 0;
        pixel_data[62][63] = 0;
        pixel_data[62][64] = 0;
        pixel_data[62][65] = 0;
        pixel_data[62][66] = 0;
        pixel_data[62][67] = 0;
        pixel_data[62][68] = 0;
        pixel_data[62][69] = 0;
        pixel_data[62][70] = 0;
        pixel_data[62][71] = 0;
        pixel_data[62][72] = 0;
        pixel_data[62][73] = 0;
        pixel_data[62][74] = 0;
        pixel_data[62][75] = 0;
        pixel_data[62][76] = 0;
        pixel_data[62][77] = 0;
        pixel_data[62][78] = 0;
        pixel_data[62][79] = 0;
        pixel_data[62][80] = 0;
        pixel_data[62][81] = 0;
        pixel_data[62][82] = 0;
        pixel_data[62][83] = 0;
        pixel_data[62][84] = 0;
        pixel_data[62][85] = 0;
        pixel_data[62][86] = 0;
        pixel_data[62][87] = 0;
        pixel_data[62][88] = 0;
        pixel_data[62][89] = 0;
        pixel_data[62][90] = 0;
        pixel_data[62][91] = 0;
        pixel_data[62][92] = 0;
        pixel_data[62][93] = 0;
        pixel_data[62][94] = 0;
        pixel_data[62][95] = 0;
        pixel_data[62][96] = 0;
        pixel_data[62][97] = 0;
        pixel_data[62][98] = 0;
        pixel_data[62][99] = 0;
        pixel_data[62][100] = 0;
        pixel_data[62][101] = 0;
        pixel_data[62][102] = 0;
        pixel_data[62][103] = 0;
        pixel_data[62][104] = 0;
        pixel_data[62][105] = 0;
        pixel_data[62][106] = 0;
        pixel_data[62][107] = 0;
        pixel_data[62][108] = 0;
        pixel_data[62][109] = 0;
        pixel_data[62][110] = 0;
        pixel_data[62][111] = 0;
        pixel_data[62][112] = 0;
        pixel_data[62][113] = 0;
        pixel_data[62][114] = 0;
        pixel_data[62][115] = 0;
        pixel_data[62][116] = 0;
        pixel_data[62][117] = 0;
        pixel_data[62][118] = 0;
        pixel_data[62][119] = 0;
        pixel_data[62][120] = 0;
        pixel_data[62][121] = 0;
        pixel_data[62][122] = 0;
        pixel_data[62][123] = 0;
        pixel_data[62][124] = 0;
        pixel_data[62][125] = 0;
        pixel_data[62][126] = 0;
        pixel_data[62][127] = 0;
        pixel_data[62][128] = 0;
        pixel_data[62][129] = 0;
        pixel_data[62][130] = 0;
        pixel_data[62][131] = 0;
        pixel_data[62][132] = 0;
        pixel_data[62][133] = 0;
        pixel_data[62][134] = 0;
        pixel_data[62][135] = 0;
        pixel_data[62][136] = 0;
        pixel_data[62][137] = 0;
        pixel_data[62][138] = 0;
        pixel_data[62][139] = 0;
        pixel_data[62][140] = 0;
        pixel_data[62][141] = 0;
        pixel_data[62][142] = 0;
        pixel_data[62][143] = 0;
        pixel_data[62][144] = 0;
        pixel_data[62][145] = 0;
        pixel_data[62][146] = 0;
        pixel_data[62][147] = 0;
        pixel_data[62][148] = 0;
        pixel_data[62][149] = 0;
        pixel_data[62][150] = 0;
        pixel_data[62][151] = 0;
        pixel_data[62][152] = 0;
        pixel_data[62][153] = 0;
        pixel_data[62][154] = 0;
        pixel_data[62][155] = 0;
        pixel_data[62][156] = 0;
        pixel_data[62][157] = 0;
        pixel_data[62][158] = 0;
        pixel_data[62][159] = 0;
        pixel_data[62][160] = 0;
        pixel_data[62][161] = 0;
        pixel_data[62][162] = 0;
        pixel_data[62][163] = 0;
        pixel_data[62][164] = 0;
        pixel_data[62][165] = 0;
        pixel_data[62][166] = 0;
        pixel_data[62][167] = 0;
        pixel_data[62][168] = 0;
        pixel_data[62][169] = 0;
        pixel_data[62][170] = 0;
        pixel_data[62][171] = 0;
        pixel_data[62][172] = 0;
        pixel_data[62][173] = 0;
        pixel_data[62][174] = 0;
        pixel_data[62][175] = 0;
        pixel_data[62][176] = 0;
        pixel_data[62][177] = 0;
        pixel_data[62][178] = 0;
        pixel_data[62][179] = 0;
        pixel_data[62][180] = 0;
        pixel_data[62][181] = 0;
        pixel_data[62][182] = 0;
        pixel_data[62][183] = 0;
        pixel_data[62][184] = 0;
        pixel_data[62][185] = 0;
        pixel_data[62][186] = 0;
        pixel_data[62][187] = 0;
        pixel_data[62][188] = 0;
        pixel_data[62][189] = 0;
        pixel_data[62][190] = 0;
        pixel_data[62][191] = 0;
        pixel_data[62][192] = 0;
        pixel_data[62][193] = 0;
        pixel_data[62][194] = 0;
        pixel_data[62][195] = 0;
        pixel_data[62][196] = 0;
        pixel_data[62][197] = 0;
        pixel_data[62][198] = 0;
        pixel_data[62][199] = 0; // y=62
        pixel_data[63][0] = 0;
        pixel_data[63][1] = 0;
        pixel_data[63][2] = 0;
        pixel_data[63][3] = 0;
        pixel_data[63][4] = 0;
        pixel_data[63][5] = 0;
        pixel_data[63][6] = 0;
        pixel_data[63][7] = 0;
        pixel_data[63][8] = 0;
        pixel_data[63][9] = 0;
        pixel_data[63][10] = 0;
        pixel_data[63][11] = 0;
        pixel_data[63][12] = 0;
        pixel_data[63][13] = 0;
        pixel_data[63][14] = 0;
        pixel_data[63][15] = 0;
        pixel_data[63][16] = 0;
        pixel_data[63][17] = 0;
        pixel_data[63][18] = 0;
        pixel_data[63][19] = 0;
        pixel_data[63][20] = 0;
        pixel_data[63][21] = 0;
        pixel_data[63][22] = 0;
        pixel_data[63][23] = 0;
        pixel_data[63][24] = 0;
        pixel_data[63][25] = 0;
        pixel_data[63][26] = 0;
        pixel_data[63][27] = 0;
        pixel_data[63][28] = 0;
        pixel_data[63][29] = 0;
        pixel_data[63][30] = 0;
        pixel_data[63][31] = 0;
        pixel_data[63][32] = 0;
        pixel_data[63][33] = 0;
        pixel_data[63][34] = 0;
        pixel_data[63][35] = 0;
        pixel_data[63][36] = 0;
        pixel_data[63][37] = 0;
        pixel_data[63][38] = 0;
        pixel_data[63][39] = 0;
        pixel_data[63][40] = 0;
        pixel_data[63][41] = 0;
        pixel_data[63][42] = 0;
        pixel_data[63][43] = 0;
        pixel_data[63][44] = 0;
        pixel_data[63][45] = 0;
        pixel_data[63][46] = 0;
        pixel_data[63][47] = 0;
        pixel_data[63][48] = 0;
        pixel_data[63][49] = 0;
        pixel_data[63][50] = 0;
        pixel_data[63][51] = 0;
        pixel_data[63][52] = 0;
        pixel_data[63][53] = 0;
        pixel_data[63][54] = 0;
        pixel_data[63][55] = 0;
        pixel_data[63][56] = 0;
        pixel_data[63][57] = 0;
        pixel_data[63][58] = 0;
        pixel_data[63][59] = 0;
        pixel_data[63][60] = 0;
        pixel_data[63][61] = 0;
        pixel_data[63][62] = 0;
        pixel_data[63][63] = 0;
        pixel_data[63][64] = 0;
        pixel_data[63][65] = 0;
        pixel_data[63][66] = 0;
        pixel_data[63][67] = 0;
        pixel_data[63][68] = 0;
        pixel_data[63][69] = 0;
        pixel_data[63][70] = 0;
        pixel_data[63][71] = 0;
        pixel_data[63][72] = 0;
        pixel_data[63][73] = 0;
        pixel_data[63][74] = 0;
        pixel_data[63][75] = 0;
        pixel_data[63][76] = 0;
        pixel_data[63][77] = 0;
        pixel_data[63][78] = 0;
        pixel_data[63][79] = 0;
        pixel_data[63][80] = 0;
        pixel_data[63][81] = 0;
        pixel_data[63][82] = 0;
        pixel_data[63][83] = 0;
        pixel_data[63][84] = 0;
        pixel_data[63][85] = 0;
        pixel_data[63][86] = 0;
        pixel_data[63][87] = 0;
        pixel_data[63][88] = 0;
        pixel_data[63][89] = 0;
        pixel_data[63][90] = 0;
        pixel_data[63][91] = 0;
        pixel_data[63][92] = 0;
        pixel_data[63][93] = 0;
        pixel_data[63][94] = 0;
        pixel_data[63][95] = 0;
        pixel_data[63][96] = 0;
        pixel_data[63][97] = 0;
        pixel_data[63][98] = 0;
        pixel_data[63][99] = 0;
        pixel_data[63][100] = 0;
        pixel_data[63][101] = 0;
        pixel_data[63][102] = 0;
        pixel_data[63][103] = 0;
        pixel_data[63][104] = 0;
        pixel_data[63][105] = 0;
        pixel_data[63][106] = 0;
        pixel_data[63][107] = 0;
        pixel_data[63][108] = 0;
        pixel_data[63][109] = 0;
        pixel_data[63][110] = 0;
        pixel_data[63][111] = 0;
        pixel_data[63][112] = 0;
        pixel_data[63][113] = 0;
        pixel_data[63][114] = 0;
        pixel_data[63][115] = 0;
        pixel_data[63][116] = 0;
        pixel_data[63][117] = 0;
        pixel_data[63][118] = 0;
        pixel_data[63][119] = 0;
        pixel_data[63][120] = 0;
        pixel_data[63][121] = 0;
        pixel_data[63][122] = 0;
        pixel_data[63][123] = 0;
        pixel_data[63][124] = 0;
        pixel_data[63][125] = 0;
        pixel_data[63][126] = 0;
        pixel_data[63][127] = 0;
        pixel_data[63][128] = 0;
        pixel_data[63][129] = 0;
        pixel_data[63][130] = 0;
        pixel_data[63][131] = 0;
        pixel_data[63][132] = 0;
        pixel_data[63][133] = 0;
        pixel_data[63][134] = 0;
        pixel_data[63][135] = 0;
        pixel_data[63][136] = 0;
        pixel_data[63][137] = 0;
        pixel_data[63][138] = 0;
        pixel_data[63][139] = 0;
        pixel_data[63][140] = 0;
        pixel_data[63][141] = 0;
        pixel_data[63][142] = 0;
        pixel_data[63][143] = 0;
        pixel_data[63][144] = 0;
        pixel_data[63][145] = 0;
        pixel_data[63][146] = 0;
        pixel_data[63][147] = 0;
        pixel_data[63][148] = 0;
        pixel_data[63][149] = 0;
        pixel_data[63][150] = 0;
        pixel_data[63][151] = 0;
        pixel_data[63][152] = 0;
        pixel_data[63][153] = 0;
        pixel_data[63][154] = 0;
        pixel_data[63][155] = 0;
        pixel_data[63][156] = 0;
        pixel_data[63][157] = 0;
        pixel_data[63][158] = 0;
        pixel_data[63][159] = 0;
        pixel_data[63][160] = 0;
        pixel_data[63][161] = 0;
        pixel_data[63][162] = 0;
        pixel_data[63][163] = 0;
        pixel_data[63][164] = 0;
        pixel_data[63][165] = 0;
        pixel_data[63][166] = 0;
        pixel_data[63][167] = 0;
        pixel_data[63][168] = 0;
        pixel_data[63][169] = 0;
        pixel_data[63][170] = 0;
        pixel_data[63][171] = 0;
        pixel_data[63][172] = 0;
        pixel_data[63][173] = 0;
        pixel_data[63][174] = 0;
        pixel_data[63][175] = 0;
        pixel_data[63][176] = 0;
        pixel_data[63][177] = 0;
        pixel_data[63][178] = 0;
        pixel_data[63][179] = 0;
        pixel_data[63][180] = 0;
        pixel_data[63][181] = 0;
        pixel_data[63][182] = 0;
        pixel_data[63][183] = 0;
        pixel_data[63][184] = 0;
        pixel_data[63][185] = 0;
        pixel_data[63][186] = 0;
        pixel_data[63][187] = 0;
        pixel_data[63][188] = 0;
        pixel_data[63][189] = 0;
        pixel_data[63][190] = 0;
        pixel_data[63][191] = 0;
        pixel_data[63][192] = 0;
        pixel_data[63][193] = 0;
        pixel_data[63][194] = 0;
        pixel_data[63][195] = 0;
        pixel_data[63][196] = 0;
        pixel_data[63][197] = 0;
        pixel_data[63][198] = 0;
        pixel_data[63][199] = 0; // y=63
        pixel_data[64][0] = 0;
        pixel_data[64][1] = 0;
        pixel_data[64][2] = 0;
        pixel_data[64][3] = 0;
        pixel_data[64][4] = 0;
        pixel_data[64][5] = 0;
        pixel_data[64][6] = 0;
        pixel_data[64][7] = 0;
        pixel_data[64][8] = 0;
        pixel_data[64][9] = 0;
        pixel_data[64][10] = 0;
        pixel_data[64][11] = 0;
        pixel_data[64][12] = 0;
        pixel_data[64][13] = 0;
        pixel_data[64][14] = 0;
        pixel_data[64][15] = 0;
        pixel_data[64][16] = 0;
        pixel_data[64][17] = 0;
        pixel_data[64][18] = 0;
        pixel_data[64][19] = 0;
        pixel_data[64][20] = 0;
        pixel_data[64][21] = 0;
        pixel_data[64][22] = 0;
        pixel_data[64][23] = 0;
        pixel_data[64][24] = 0;
        pixel_data[64][25] = 0;
        pixel_data[64][26] = 0;
        pixel_data[64][27] = 0;
        pixel_data[64][28] = 0;
        pixel_data[64][29] = 0;
        pixel_data[64][30] = 0;
        pixel_data[64][31] = 0;
        pixel_data[64][32] = 0;
        pixel_data[64][33] = 0;
        pixel_data[64][34] = 0;
        pixel_data[64][35] = 0;
        pixel_data[64][36] = 0;
        pixel_data[64][37] = 0;
        pixel_data[64][38] = 0;
        pixel_data[64][39] = 0;
        pixel_data[64][40] = 0;
        pixel_data[64][41] = 0;
        pixel_data[64][42] = 0;
        pixel_data[64][43] = 0;
        pixel_data[64][44] = 0;
        pixel_data[64][45] = 0;
        pixel_data[64][46] = 0;
        pixel_data[64][47] = 0;
        pixel_data[64][48] = 0;
        pixel_data[64][49] = 0;
        pixel_data[64][50] = 0;
        pixel_data[64][51] = 0;
        pixel_data[64][52] = 0;
        pixel_data[64][53] = 0;
        pixel_data[64][54] = 0;
        pixel_data[64][55] = 0;
        pixel_data[64][56] = 0;
        pixel_data[64][57] = 0;
        pixel_data[64][58] = 0;
        pixel_data[64][59] = 0;
        pixel_data[64][60] = 0;
        pixel_data[64][61] = 0;
        pixel_data[64][62] = 0;
        pixel_data[64][63] = 0;
        pixel_data[64][64] = 0;
        pixel_data[64][65] = 0;
        pixel_data[64][66] = 0;
        pixel_data[64][67] = 0;
        pixel_data[64][68] = 0;
        pixel_data[64][69] = 0;
        pixel_data[64][70] = 0;
        pixel_data[64][71] = 0;
        pixel_data[64][72] = 0;
        pixel_data[64][73] = 0;
        pixel_data[64][74] = 0;
        pixel_data[64][75] = 0;
        pixel_data[64][76] = 0;
        pixel_data[64][77] = 0;
        pixel_data[64][78] = 0;
        pixel_data[64][79] = 0;
        pixel_data[64][80] = 0;
        pixel_data[64][81] = 0;
        pixel_data[64][82] = 0;
        pixel_data[64][83] = 0;
        pixel_data[64][84] = 0;
        pixel_data[64][85] = 0;
        pixel_data[64][86] = 0;
        pixel_data[64][87] = 0;
        pixel_data[64][88] = 0;
        pixel_data[64][89] = 0;
        pixel_data[64][90] = 0;
        pixel_data[64][91] = 0;
        pixel_data[64][92] = 0;
        pixel_data[64][93] = 0;
        pixel_data[64][94] = 0;
        pixel_data[64][95] = 0;
        pixel_data[64][96] = 0;
        pixel_data[64][97] = 0;
        pixel_data[64][98] = 0;
        pixel_data[64][99] = 0;
        pixel_data[64][100] = 0;
        pixel_data[64][101] = 0;
        pixel_data[64][102] = 0;
        pixel_data[64][103] = 0;
        pixel_data[64][104] = 0;
        pixel_data[64][105] = 0;
        pixel_data[64][106] = 0;
        pixel_data[64][107] = 0;
        pixel_data[64][108] = 0;
        pixel_data[64][109] = 0;
        pixel_data[64][110] = 0;
        pixel_data[64][111] = 0;
        pixel_data[64][112] = 0;
        pixel_data[64][113] = 0;
        pixel_data[64][114] = 0;
        pixel_data[64][115] = 0;
        pixel_data[64][116] = 0;
        pixel_data[64][117] = 0;
        pixel_data[64][118] = 0;
        pixel_data[64][119] = 0;
        pixel_data[64][120] = 0;
        pixel_data[64][121] = 0;
        pixel_data[64][122] = 0;
        pixel_data[64][123] = 0;
        pixel_data[64][124] = 0;
        pixel_data[64][125] = 0;
        pixel_data[64][126] = 0;
        pixel_data[64][127] = 0;
        pixel_data[64][128] = 0;
        pixel_data[64][129] = 0;
        pixel_data[64][130] = 0;
        pixel_data[64][131] = 0;
        pixel_data[64][132] = 0;
        pixel_data[64][133] = 0;
        pixel_data[64][134] = 0;
        pixel_data[64][135] = 0;
        pixel_data[64][136] = 0;
        pixel_data[64][137] = 0;
        pixel_data[64][138] = 0;
        pixel_data[64][139] = 0;
        pixel_data[64][140] = 0;
        pixel_data[64][141] = 0;
        pixel_data[64][142] = 0;
        pixel_data[64][143] = 0;
        pixel_data[64][144] = 0;
        pixel_data[64][145] = 0;
        pixel_data[64][146] = 0;
        pixel_data[64][147] = 0;
        pixel_data[64][148] = 0;
        pixel_data[64][149] = 0;
        pixel_data[64][150] = 0;
        pixel_data[64][151] = 0;
        pixel_data[64][152] = 0;
        pixel_data[64][153] = 0;
        pixel_data[64][154] = 0;
        pixel_data[64][155] = 0;
        pixel_data[64][156] = 0;
        pixel_data[64][157] = 0;
        pixel_data[64][158] = 0;
        pixel_data[64][159] = 0;
        pixel_data[64][160] = 0;
        pixel_data[64][161] = 0;
        pixel_data[64][162] = 0;
        pixel_data[64][163] = 0;
        pixel_data[64][164] = 0;
        pixel_data[64][165] = 0;
        pixel_data[64][166] = 0;
        pixel_data[64][167] = 0;
        pixel_data[64][168] = 0;
        pixel_data[64][169] = 0;
        pixel_data[64][170] = 0;
        pixel_data[64][171] = 0;
        pixel_data[64][172] = 0;
        pixel_data[64][173] = 0;
        pixel_data[64][174] = 0;
        pixel_data[64][175] = 0;
        pixel_data[64][176] = 0;
        pixel_data[64][177] = 0;
        pixel_data[64][178] = 0;
        pixel_data[64][179] = 0;
        pixel_data[64][180] = 0;
        pixel_data[64][181] = 0;
        pixel_data[64][182] = 0;
        pixel_data[64][183] = 0;
        pixel_data[64][184] = 0;
        pixel_data[64][185] = 0;
        pixel_data[64][186] = 0;
        pixel_data[64][187] = 0;
        pixel_data[64][188] = 0;
        pixel_data[64][189] = 0;
        pixel_data[64][190] = 0;
        pixel_data[64][191] = 0;
        pixel_data[64][192] = 0;
        pixel_data[64][193] = 0;
        pixel_data[64][194] = 0;
        pixel_data[64][195] = 0;
        pixel_data[64][196] = 0;
        pixel_data[64][197] = 0;
        pixel_data[64][198] = 0;
        pixel_data[64][199] = 0; // y=64
        pixel_data[65][0] = 0;
        pixel_data[65][1] = 0;
        pixel_data[65][2] = 0;
        pixel_data[65][3] = 0;
        pixel_data[65][4] = 0;
        pixel_data[65][5] = 0;
        pixel_data[65][6] = 0;
        pixel_data[65][7] = 0;
        pixel_data[65][8] = 0;
        pixel_data[65][9] = 0;
        pixel_data[65][10] = 0;
        pixel_data[65][11] = 0;
        pixel_data[65][12] = 0;
        pixel_data[65][13] = 0;
        pixel_data[65][14] = 0;
        pixel_data[65][15] = 0;
        pixel_data[65][16] = 0;
        pixel_data[65][17] = 0;
        pixel_data[65][18] = 0;
        pixel_data[65][19] = 0;
        pixel_data[65][20] = 0;
        pixel_data[65][21] = 0;
        pixel_data[65][22] = 0;
        pixel_data[65][23] = 0;
        pixel_data[65][24] = 0;
        pixel_data[65][25] = 0;
        pixel_data[65][26] = 0;
        pixel_data[65][27] = 0;
        pixel_data[65][28] = 0;
        pixel_data[65][29] = 0;
        pixel_data[65][30] = 0;
        pixel_data[65][31] = 0;
        pixel_data[65][32] = 0;
        pixel_data[65][33] = 0;
        pixel_data[65][34] = 0;
        pixel_data[65][35] = 0;
        pixel_data[65][36] = 0;
        pixel_data[65][37] = 0;
        pixel_data[65][38] = 0;
        pixel_data[65][39] = 0;
        pixel_data[65][40] = 0;
        pixel_data[65][41] = 0;
        pixel_data[65][42] = 0;
        pixel_data[65][43] = 0;
        pixel_data[65][44] = 0;
        pixel_data[65][45] = 0;
        pixel_data[65][46] = 0;
        pixel_data[65][47] = 0;
        pixel_data[65][48] = 0;
        pixel_data[65][49] = 0;
        pixel_data[65][50] = 0;
        pixel_data[65][51] = 0;
        pixel_data[65][52] = 0;
        pixel_data[65][53] = 0;
        pixel_data[65][54] = 0;
        pixel_data[65][55] = 0;
        pixel_data[65][56] = 0;
        pixel_data[65][57] = 0;
        pixel_data[65][58] = 0;
        pixel_data[65][59] = 0;
        pixel_data[65][60] = 0;
        pixel_data[65][61] = 0;
        pixel_data[65][62] = 0;
        pixel_data[65][63] = 0;
        pixel_data[65][64] = 0;
        pixel_data[65][65] = 0;
        pixel_data[65][66] = 0;
        pixel_data[65][67] = 0;
        pixel_data[65][68] = 0;
        pixel_data[65][69] = 0;
        pixel_data[65][70] = 0;
        pixel_data[65][71] = 0;
        pixel_data[65][72] = 0;
        pixel_data[65][73] = 0;
        pixel_data[65][74] = 0;
        pixel_data[65][75] = 0;
        pixel_data[65][76] = 0;
        pixel_data[65][77] = 0;
        pixel_data[65][78] = 0;
        pixel_data[65][79] = 0;
        pixel_data[65][80] = 0;
        pixel_data[65][81] = 0;
        pixel_data[65][82] = 0;
        pixel_data[65][83] = 0;
        pixel_data[65][84] = 0;
        pixel_data[65][85] = 0;
        pixel_data[65][86] = 0;
        pixel_data[65][87] = 0;
        pixel_data[65][88] = 0;
        pixel_data[65][89] = 0;
        pixel_data[65][90] = 0;
        pixel_data[65][91] = 0;
        pixel_data[65][92] = 0;
        pixel_data[65][93] = 0;
        pixel_data[65][94] = 0;
        pixel_data[65][95] = 0;
        pixel_data[65][96] = 0;
        pixel_data[65][97] = 0;
        pixel_data[65][98] = 0;
        pixel_data[65][99] = 0;
        pixel_data[65][100] = 0;
        pixel_data[65][101] = 0;
        pixel_data[65][102] = 0;
        pixel_data[65][103] = 0;
        pixel_data[65][104] = 0;
        pixel_data[65][105] = 0;
        pixel_data[65][106] = 0;
        pixel_data[65][107] = 0;
        pixel_data[65][108] = 0;
        pixel_data[65][109] = 0;
        pixel_data[65][110] = 0;
        pixel_data[65][111] = 0;
        pixel_data[65][112] = 0;
        pixel_data[65][113] = 0;
        pixel_data[65][114] = 0;
        pixel_data[65][115] = 0;
        pixel_data[65][116] = 0;
        pixel_data[65][117] = 0;
        pixel_data[65][118] = 0;
        pixel_data[65][119] = 0;
        pixel_data[65][120] = 0;
        pixel_data[65][121] = 0;
        pixel_data[65][122] = 0;
        pixel_data[65][123] = 0;
        pixel_data[65][124] = 0;
        pixel_data[65][125] = 0;
        pixel_data[65][126] = 0;
        pixel_data[65][127] = 0;
        pixel_data[65][128] = 0;
        pixel_data[65][129] = 0;
        pixel_data[65][130] = 0;
        pixel_data[65][131] = 0;
        pixel_data[65][132] = 0;
        pixel_data[65][133] = 0;
        pixel_data[65][134] = 0;
        pixel_data[65][135] = 0;
        pixel_data[65][136] = 0;
        pixel_data[65][137] = 0;
        pixel_data[65][138] = 0;
        pixel_data[65][139] = 0;
        pixel_data[65][140] = 0;
        pixel_data[65][141] = 0;
        pixel_data[65][142] = 0;
        pixel_data[65][143] = 0;
        pixel_data[65][144] = 0;
        pixel_data[65][145] = 0;
        pixel_data[65][146] = 0;
        pixel_data[65][147] = 0;
        pixel_data[65][148] = 0;
        pixel_data[65][149] = 0;
        pixel_data[65][150] = 0;
        pixel_data[65][151] = 0;
        pixel_data[65][152] = 0;
        pixel_data[65][153] = 0;
        pixel_data[65][154] = 0;
        pixel_data[65][155] = 0;
        pixel_data[65][156] = 0;
        pixel_data[65][157] = 0;
        pixel_data[65][158] = 0;
        pixel_data[65][159] = 0;
        pixel_data[65][160] = 0;
        pixel_data[65][161] = 0;
        pixel_data[65][162] = 0;
        pixel_data[65][163] = 0;
        pixel_data[65][164] = 0;
        pixel_data[65][165] = 0;
        pixel_data[65][166] = 0;
        pixel_data[65][167] = 0;
        pixel_data[65][168] = 0;
        pixel_data[65][169] = 0;
        pixel_data[65][170] = 0;
        pixel_data[65][171] = 0;
        pixel_data[65][172] = 0;
        pixel_data[65][173] = 0;
        pixel_data[65][174] = 0;
        pixel_data[65][175] = 0;
        pixel_data[65][176] = 0;
        pixel_data[65][177] = 0;
        pixel_data[65][178] = 0;
        pixel_data[65][179] = 0;
        pixel_data[65][180] = 0;
        pixel_data[65][181] = 0;
        pixel_data[65][182] = 0;
        pixel_data[65][183] = 0;
        pixel_data[65][184] = 0;
        pixel_data[65][185] = 0;
        pixel_data[65][186] = 0;
        pixel_data[65][187] = 0;
        pixel_data[65][188] = 0;
        pixel_data[65][189] = 0;
        pixel_data[65][190] = 0;
        pixel_data[65][191] = 0;
        pixel_data[65][192] = 0;
        pixel_data[65][193] = 0;
        pixel_data[65][194] = 0;
        pixel_data[65][195] = 0;
        pixel_data[65][196] = 0;
        pixel_data[65][197] = 0;
        pixel_data[65][198] = 0;
        pixel_data[65][199] = 0; // y=65
        pixel_data[66][0] = 0;
        pixel_data[66][1] = 0;
        pixel_data[66][2] = 0;
        pixel_data[66][3] = 0;
        pixel_data[66][4] = 0;
        pixel_data[66][5] = 0;
        pixel_data[66][6] = 0;
        pixel_data[66][7] = 0;
        pixel_data[66][8] = 0;
        pixel_data[66][9] = 0;
        pixel_data[66][10] = 0;
        pixel_data[66][11] = 0;
        pixel_data[66][12] = 0;
        pixel_data[66][13] = 0;
        pixel_data[66][14] = 0;
        pixel_data[66][15] = 0;
        pixel_data[66][16] = 0;
        pixel_data[66][17] = 0;
        pixel_data[66][18] = 0;
        pixel_data[66][19] = 0;
        pixel_data[66][20] = 0;
        pixel_data[66][21] = 0;
        pixel_data[66][22] = 0;
        pixel_data[66][23] = 0;
        pixel_data[66][24] = 0;
        pixel_data[66][25] = 0;
        pixel_data[66][26] = 0;
        pixel_data[66][27] = 0;
        pixel_data[66][28] = 0;
        pixel_data[66][29] = 0;
        pixel_data[66][30] = 0;
        pixel_data[66][31] = 0;
        pixel_data[66][32] = 0;
        pixel_data[66][33] = 0;
        pixel_data[66][34] = 0;
        pixel_data[66][35] = 0;
        pixel_data[66][36] = 0;
        pixel_data[66][37] = 0;
        pixel_data[66][38] = 0;
        pixel_data[66][39] = 0;
        pixel_data[66][40] = 0;
        pixel_data[66][41] = 0;
        pixel_data[66][42] = 0;
        pixel_data[66][43] = 0;
        pixel_data[66][44] = 0;
        pixel_data[66][45] = 0;
        pixel_data[66][46] = 0;
        pixel_data[66][47] = 0;
        pixel_data[66][48] = 0;
        pixel_data[66][49] = 0;
        pixel_data[66][50] = 0;
        pixel_data[66][51] = 0;
        pixel_data[66][52] = 0;
        pixel_data[66][53] = 0;
        pixel_data[66][54] = 0;
        pixel_data[66][55] = 0;
        pixel_data[66][56] = 0;
        pixel_data[66][57] = 0;
        pixel_data[66][58] = 0;
        pixel_data[66][59] = 0;
        pixel_data[66][60] = 0;
        pixel_data[66][61] = 0;
        pixel_data[66][62] = 0;
        pixel_data[66][63] = 0;
        pixel_data[66][64] = 0;
        pixel_data[66][65] = 0;
        pixel_data[66][66] = 0;
        pixel_data[66][67] = 0;
        pixel_data[66][68] = 0;
        pixel_data[66][69] = 0;
        pixel_data[66][70] = 0;
        pixel_data[66][71] = 0;
        pixel_data[66][72] = 0;
        pixel_data[66][73] = 0;
        pixel_data[66][74] = 0;
        pixel_data[66][75] = 0;
        pixel_data[66][76] = 0;
        pixel_data[66][77] = 0;
        pixel_data[66][78] = 0;
        pixel_data[66][79] = 0;
        pixel_data[66][80] = 0;
        pixel_data[66][81] = 0;
        pixel_data[66][82] = 0;
        pixel_data[66][83] = 0;
        pixel_data[66][84] = 0;
        pixel_data[66][85] = 0;
        pixel_data[66][86] = 0;
        pixel_data[66][87] = 0;
        pixel_data[66][88] = 0;
        pixel_data[66][89] = 0;
        pixel_data[66][90] = 0;
        pixel_data[66][91] = 0;
        pixel_data[66][92] = 0;
        pixel_data[66][93] = 0;
        pixel_data[66][94] = 0;
        pixel_data[66][95] = 0;
        pixel_data[66][96] = 0;
        pixel_data[66][97] = 0;
        pixel_data[66][98] = 0;
        pixel_data[66][99] = 0;
        pixel_data[66][100] = 0;
        pixel_data[66][101] = 0;
        pixel_data[66][102] = 0;
        pixel_data[66][103] = 0;
        pixel_data[66][104] = 0;
        pixel_data[66][105] = 0;
        pixel_data[66][106] = 0;
        pixel_data[66][107] = 0;
        pixel_data[66][108] = 0;
        pixel_data[66][109] = 0;
        pixel_data[66][110] = 0;
        pixel_data[66][111] = 0;
        pixel_data[66][112] = 0;
        pixel_data[66][113] = 0;
        pixel_data[66][114] = 0;
        pixel_data[66][115] = 0;
        pixel_data[66][116] = 0;
        pixel_data[66][117] = 0;
        pixel_data[66][118] = 0;
        pixel_data[66][119] = 0;
        pixel_data[66][120] = 0;
        pixel_data[66][121] = 0;
        pixel_data[66][122] = 0;
        pixel_data[66][123] = 0;
        pixel_data[66][124] = 0;
        pixel_data[66][125] = 0;
        pixel_data[66][126] = 0;
        pixel_data[66][127] = 0;
        pixel_data[66][128] = 0;
        pixel_data[66][129] = 0;
        pixel_data[66][130] = 0;
        pixel_data[66][131] = 0;
        pixel_data[66][132] = 0;
        pixel_data[66][133] = 0;
        pixel_data[66][134] = 0;
        pixel_data[66][135] = 0;
        pixel_data[66][136] = 0;
        pixel_data[66][137] = 0;
        pixel_data[66][138] = 0;
        pixel_data[66][139] = 0;
        pixel_data[66][140] = 0;
        pixel_data[66][141] = 0;
        pixel_data[66][142] = 0;
        pixel_data[66][143] = 0;
        pixel_data[66][144] = 0;
        pixel_data[66][145] = 0;
        pixel_data[66][146] = 0;
        pixel_data[66][147] = 0;
        pixel_data[66][148] = 0;
        pixel_data[66][149] = 0;
        pixel_data[66][150] = 0;
        pixel_data[66][151] = 0;
        pixel_data[66][152] = 0;
        pixel_data[66][153] = 0;
        pixel_data[66][154] = 0;
        pixel_data[66][155] = 0;
        pixel_data[66][156] = 0;
        pixel_data[66][157] = 0;
        pixel_data[66][158] = 0;
        pixel_data[66][159] = 0;
        pixel_data[66][160] = 0;
        pixel_data[66][161] = 0;
        pixel_data[66][162] = 0;
        pixel_data[66][163] = 0;
        pixel_data[66][164] = 0;
        pixel_data[66][165] = 0;
        pixel_data[66][166] = 0;
        pixel_data[66][167] = 0;
        pixel_data[66][168] = 0;
        pixel_data[66][169] = 0;
        pixel_data[66][170] = 0;
        pixel_data[66][171] = 0;
        pixel_data[66][172] = 0;
        pixel_data[66][173] = 0;
        pixel_data[66][174] = 0;
        pixel_data[66][175] = 0;
        pixel_data[66][176] = 0;
        pixel_data[66][177] = 0;
        pixel_data[66][178] = 0;
        pixel_data[66][179] = 0;
        pixel_data[66][180] = 0;
        pixel_data[66][181] = 0;
        pixel_data[66][182] = 0;
        pixel_data[66][183] = 0;
        pixel_data[66][184] = 0;
        pixel_data[66][185] = 0;
        pixel_data[66][186] = 0;
        pixel_data[66][187] = 0;
        pixel_data[66][188] = 0;
        pixel_data[66][189] = 0;
        pixel_data[66][190] = 0;
        pixel_data[66][191] = 0;
        pixel_data[66][192] = 0;
        pixel_data[66][193] = 0;
        pixel_data[66][194] = 0;
        pixel_data[66][195] = 0;
        pixel_data[66][196] = 0;
        pixel_data[66][197] = 0;
        pixel_data[66][198] = 0;
        pixel_data[66][199] = 0; // y=66
        pixel_data[67][0] = 0;
        pixel_data[67][1] = 0;
        pixel_data[67][2] = 0;
        pixel_data[67][3] = 0;
        pixel_data[67][4] = 0;
        pixel_data[67][5] = 0;
        pixel_data[67][6] = 0;
        pixel_data[67][7] = 0;
        pixel_data[67][8] = 0;
        pixel_data[67][9] = 0;
        pixel_data[67][10] = 0;
        pixel_data[67][11] = 0;
        pixel_data[67][12] = 0;
        pixel_data[67][13] = 0;
        pixel_data[67][14] = 0;
        pixel_data[67][15] = 0;
        pixel_data[67][16] = 0;
        pixel_data[67][17] = 0;
        pixel_data[67][18] = 0;
        pixel_data[67][19] = 0;
        pixel_data[67][20] = 0;
        pixel_data[67][21] = 0;
        pixel_data[67][22] = 0;
        pixel_data[67][23] = 0;
        pixel_data[67][24] = 0;
        pixel_data[67][25] = 0;
        pixel_data[67][26] = 0;
        pixel_data[67][27] = 0;
        pixel_data[67][28] = 0;
        pixel_data[67][29] = 0;
        pixel_data[67][30] = 0;
        pixel_data[67][31] = 0;
        pixel_data[67][32] = 0;
        pixel_data[67][33] = 0;
        pixel_data[67][34] = 0;
        pixel_data[67][35] = 0;
        pixel_data[67][36] = 0;
        pixel_data[67][37] = 0;
        pixel_data[67][38] = 0;
        pixel_data[67][39] = 0;
        pixel_data[67][40] = 0;
        pixel_data[67][41] = 0;
        pixel_data[67][42] = 0;
        pixel_data[67][43] = 0;
        pixel_data[67][44] = 0;
        pixel_data[67][45] = 0;
        pixel_data[67][46] = 0;
        pixel_data[67][47] = 0;
        pixel_data[67][48] = 0;
        pixel_data[67][49] = 0;
        pixel_data[67][50] = 0;
        pixel_data[67][51] = 0;
        pixel_data[67][52] = 0;
        pixel_data[67][53] = 0;
        pixel_data[67][54] = 0;
        pixel_data[67][55] = 0;
        pixel_data[67][56] = 0;
        pixel_data[67][57] = 0;
        pixel_data[67][58] = 0;
        pixel_data[67][59] = 0;
        pixel_data[67][60] = 0;
        pixel_data[67][61] = 0;
        pixel_data[67][62] = 0;
        pixel_data[67][63] = 0;
        pixel_data[67][64] = 0;
        pixel_data[67][65] = 0;
        pixel_data[67][66] = 0;
        pixel_data[67][67] = 0;
        pixel_data[67][68] = 0;
        pixel_data[67][69] = 0;
        pixel_data[67][70] = 0;
        pixel_data[67][71] = 0;
        pixel_data[67][72] = 0;
        pixel_data[67][73] = 0;
        pixel_data[67][74] = 0;
        pixel_data[67][75] = 0;
        pixel_data[67][76] = 0;
        pixel_data[67][77] = 0;
        pixel_data[67][78] = 0;
        pixel_data[67][79] = 0;
        pixel_data[67][80] = 0;
        pixel_data[67][81] = 0;
        pixel_data[67][82] = 0;
        pixel_data[67][83] = 0;
        pixel_data[67][84] = 0;
        pixel_data[67][85] = 0;
        pixel_data[67][86] = 0;
        pixel_data[67][87] = 0;
        pixel_data[67][88] = 0;
        pixel_data[67][89] = 0;
        pixel_data[67][90] = 0;
        pixel_data[67][91] = 0;
        pixel_data[67][92] = 0;
        pixel_data[67][93] = 0;
        pixel_data[67][94] = 0;
        pixel_data[67][95] = 0;
        pixel_data[67][96] = 0;
        pixel_data[67][97] = 0;
        pixel_data[67][98] = 0;
        pixel_data[67][99] = 0;
        pixel_data[67][100] = 0;
        pixel_data[67][101] = 0;
        pixel_data[67][102] = 0;
        pixel_data[67][103] = 0;
        pixel_data[67][104] = 0;
        pixel_data[67][105] = 0;
        pixel_data[67][106] = 0;
        pixel_data[67][107] = 0;
        pixel_data[67][108] = 0;
        pixel_data[67][109] = 0;
        pixel_data[67][110] = 0;
        pixel_data[67][111] = 0;
        pixel_data[67][112] = 0;
        pixel_data[67][113] = 0;
        pixel_data[67][114] = 0;
        pixel_data[67][115] = 0;
        pixel_data[67][116] = 0;
        pixel_data[67][117] = 0;
        pixel_data[67][118] = 0;
        pixel_data[67][119] = 0;
        pixel_data[67][120] = 0;
        pixel_data[67][121] = 0;
        pixel_data[67][122] = 0;
        pixel_data[67][123] = 0;
        pixel_data[67][124] = 0;
        pixel_data[67][125] = 0;
        pixel_data[67][126] = 0;
        pixel_data[67][127] = 0;
        pixel_data[67][128] = 0;
        pixel_data[67][129] = 0;
        pixel_data[67][130] = 0;
        pixel_data[67][131] = 0;
        pixel_data[67][132] = 0;
        pixel_data[67][133] = 0;
        pixel_data[67][134] = 0;
        pixel_data[67][135] = 0;
        pixel_data[67][136] = 0;
        pixel_data[67][137] = 0;
        pixel_data[67][138] = 0;
        pixel_data[67][139] = 0;
        pixel_data[67][140] = 0;
        pixel_data[67][141] = 0;
        pixel_data[67][142] = 0;
        pixel_data[67][143] = 0;
        pixel_data[67][144] = 0;
        pixel_data[67][145] = 0;
        pixel_data[67][146] = 0;
        pixel_data[67][147] = 0;
        pixel_data[67][148] = 0;
        pixel_data[67][149] = 0;
        pixel_data[67][150] = 0;
        pixel_data[67][151] = 0;
        pixel_data[67][152] = 0;
        pixel_data[67][153] = 0;
        pixel_data[67][154] = 0;
        pixel_data[67][155] = 0;
        pixel_data[67][156] = 0;
        pixel_data[67][157] = 0;
        pixel_data[67][158] = 0;
        pixel_data[67][159] = 0;
        pixel_data[67][160] = 0;
        pixel_data[67][161] = 0;
        pixel_data[67][162] = 0;
        pixel_data[67][163] = 0;
        pixel_data[67][164] = 0;
        pixel_data[67][165] = 0;
        pixel_data[67][166] = 0;
        pixel_data[67][167] = 0;
        pixel_data[67][168] = 0;
        pixel_data[67][169] = 0;
        pixel_data[67][170] = 0;
        pixel_data[67][171] = 0;
        pixel_data[67][172] = 0;
        pixel_data[67][173] = 0;
        pixel_data[67][174] = 0;
        pixel_data[67][175] = 0;
        pixel_data[67][176] = 0;
        pixel_data[67][177] = 0;
        pixel_data[67][178] = 0;
        pixel_data[67][179] = 0;
        pixel_data[67][180] = 0;
        pixel_data[67][181] = 0;
        pixel_data[67][182] = 0;
        pixel_data[67][183] = 0;
        pixel_data[67][184] = 0;
        pixel_data[67][185] = 0;
        pixel_data[67][186] = 0;
        pixel_data[67][187] = 0;
        pixel_data[67][188] = 0;
        pixel_data[67][189] = 0;
        pixel_data[67][190] = 0;
        pixel_data[67][191] = 0;
        pixel_data[67][192] = 0;
        pixel_data[67][193] = 0;
        pixel_data[67][194] = 0;
        pixel_data[67][195] = 0;
        pixel_data[67][196] = 0;
        pixel_data[67][197] = 0;
        pixel_data[67][198] = 0;
        pixel_data[67][199] = 0; // y=67
        pixel_data[68][0] = 0;
        pixel_data[68][1] = 0;
        pixel_data[68][2] = 0;
        pixel_data[68][3] = 0;
        pixel_data[68][4] = 0;
        pixel_data[68][5] = 0;
        pixel_data[68][6] = 0;
        pixel_data[68][7] = 0;
        pixel_data[68][8] = 0;
        pixel_data[68][9] = 0;
        pixel_data[68][10] = 0;
        pixel_data[68][11] = 0;
        pixel_data[68][12] = 0;
        pixel_data[68][13] = 0;
        pixel_data[68][14] = 0;
        pixel_data[68][15] = 0;
        pixel_data[68][16] = 0;
        pixel_data[68][17] = 0;
        pixel_data[68][18] = 0;
        pixel_data[68][19] = 0;
        pixel_data[68][20] = 0;
        pixel_data[68][21] = 0;
        pixel_data[68][22] = 0;
        pixel_data[68][23] = 0;
        pixel_data[68][24] = 0;
        pixel_data[68][25] = 0;
        pixel_data[68][26] = 0;
        pixel_data[68][27] = 0;
        pixel_data[68][28] = 0;
        pixel_data[68][29] = 0;
        pixel_data[68][30] = 0;
        pixel_data[68][31] = 0;
        pixel_data[68][32] = 0;
        pixel_data[68][33] = 0;
        pixel_data[68][34] = 0;
        pixel_data[68][35] = 0;
        pixel_data[68][36] = 0;
        pixel_data[68][37] = 0;
        pixel_data[68][38] = 0;
        pixel_data[68][39] = 0;
        pixel_data[68][40] = 0;
        pixel_data[68][41] = 0;
        pixel_data[68][42] = 0;
        pixel_data[68][43] = 0;
        pixel_data[68][44] = 0;
        pixel_data[68][45] = 0;
        pixel_data[68][46] = 0;
        pixel_data[68][47] = 0;
        pixel_data[68][48] = 0;
        pixel_data[68][49] = 0;
        pixel_data[68][50] = 0;
        pixel_data[68][51] = 0;
        pixel_data[68][52] = 0;
        pixel_data[68][53] = 0;
        pixel_data[68][54] = 0;
        pixel_data[68][55] = 0;
        pixel_data[68][56] = 0;
        pixel_data[68][57] = 0;
        pixel_data[68][58] = 0;
        pixel_data[68][59] = 0;
        pixel_data[68][60] = 0;
        pixel_data[68][61] = 0;
        pixel_data[68][62] = 0;
        pixel_data[68][63] = 0;
        pixel_data[68][64] = 0;
        pixel_data[68][65] = 0;
        pixel_data[68][66] = 0;
        pixel_data[68][67] = 0;
        pixel_data[68][68] = 0;
        pixel_data[68][69] = 0;
        pixel_data[68][70] = 0;
        pixel_data[68][71] = 0;
        pixel_data[68][72] = 0;
        pixel_data[68][73] = 0;
        pixel_data[68][74] = 0;
        pixel_data[68][75] = 0;
        pixel_data[68][76] = 0;
        pixel_data[68][77] = 0;
        pixel_data[68][78] = 0;
        pixel_data[68][79] = 0;
        pixel_data[68][80] = 0;
        pixel_data[68][81] = 0;
        pixel_data[68][82] = 0;
        pixel_data[68][83] = 0;
        pixel_data[68][84] = 0;
        pixel_data[68][85] = 0;
        pixel_data[68][86] = 0;
        pixel_data[68][87] = 0;
        pixel_data[68][88] = 0;
        pixel_data[68][89] = 0;
        pixel_data[68][90] = 0;
        pixel_data[68][91] = 0;
        pixel_data[68][92] = 0;
        pixel_data[68][93] = 0;
        pixel_data[68][94] = 0;
        pixel_data[68][95] = 0;
        pixel_data[68][96] = 0;
        pixel_data[68][97] = 0;
        pixel_data[68][98] = 0;
        pixel_data[68][99] = 0;
        pixel_data[68][100] = 0;
        pixel_data[68][101] = 0;
        pixel_data[68][102] = 0;
        pixel_data[68][103] = 0;
        pixel_data[68][104] = 0;
        pixel_data[68][105] = 0;
        pixel_data[68][106] = 0;
        pixel_data[68][107] = 0;
        pixel_data[68][108] = 0;
        pixel_data[68][109] = 0;
        pixel_data[68][110] = 0;
        pixel_data[68][111] = 0;
        pixel_data[68][112] = 0;
        pixel_data[68][113] = 0;
        pixel_data[68][114] = 0;
        pixel_data[68][115] = 0;
        pixel_data[68][116] = 0;
        pixel_data[68][117] = 0;
        pixel_data[68][118] = 0;
        pixel_data[68][119] = 0;
        pixel_data[68][120] = 0;
        pixel_data[68][121] = 0;
        pixel_data[68][122] = 0;
        pixel_data[68][123] = 0;
        pixel_data[68][124] = 0;
        pixel_data[68][125] = 0;
        pixel_data[68][126] = 0;
        pixel_data[68][127] = 0;
        pixel_data[68][128] = 0;
        pixel_data[68][129] = 0;
        pixel_data[68][130] = 0;
        pixel_data[68][131] = 0;
        pixel_data[68][132] = 0;
        pixel_data[68][133] = 0;
        pixel_data[68][134] = 0;
        pixel_data[68][135] = 0;
        pixel_data[68][136] = 0;
        pixel_data[68][137] = 0;
        pixel_data[68][138] = 0;
        pixel_data[68][139] = 0;
        pixel_data[68][140] = 0;
        pixel_data[68][141] = 0;
        pixel_data[68][142] = 0;
        pixel_data[68][143] = 0;
        pixel_data[68][144] = 0;
        pixel_data[68][145] = 0;
        pixel_data[68][146] = 0;
        pixel_data[68][147] = 0;
        pixel_data[68][148] = 0;
        pixel_data[68][149] = 0;
        pixel_data[68][150] = 0;
        pixel_data[68][151] = 0;
        pixel_data[68][152] = 0;
        pixel_data[68][153] = 0;
        pixel_data[68][154] = 0;
        pixel_data[68][155] = 0;
        pixel_data[68][156] = 0;
        pixel_data[68][157] = 0;
        pixel_data[68][158] = 0;
        pixel_data[68][159] = 0;
        pixel_data[68][160] = 0;
        pixel_data[68][161] = 0;
        pixel_data[68][162] = 0;
        pixel_data[68][163] = 0;
        pixel_data[68][164] = 0;
        pixel_data[68][165] = 0;
        pixel_data[68][166] = 0;
        pixel_data[68][167] = 0;
        pixel_data[68][168] = 0;
        pixel_data[68][169] = 0;
        pixel_data[68][170] = 0;
        pixel_data[68][171] = 0;
        pixel_data[68][172] = 0;
        pixel_data[68][173] = 0;
        pixel_data[68][174] = 0;
        pixel_data[68][175] = 0;
        pixel_data[68][176] = 0;
        pixel_data[68][177] = 0;
        pixel_data[68][178] = 0;
        pixel_data[68][179] = 0;
        pixel_data[68][180] = 0;
        pixel_data[68][181] = 0;
        pixel_data[68][182] = 0;
        pixel_data[68][183] = 0;
        pixel_data[68][184] = 0;
        pixel_data[68][185] = 0;
        pixel_data[68][186] = 0;
        pixel_data[68][187] = 0;
        pixel_data[68][188] = 0;
        pixel_data[68][189] = 0;
        pixel_data[68][190] = 0;
        pixel_data[68][191] = 0;
        pixel_data[68][192] = 0;
        pixel_data[68][193] = 0;
        pixel_data[68][194] = 0;
        pixel_data[68][195] = 0;
        pixel_data[68][196] = 0;
        pixel_data[68][197] = 0;
        pixel_data[68][198] = 0;
        pixel_data[68][199] = 0; // y=68
        pixel_data[69][0] = 0;
        pixel_data[69][1] = 0;
        pixel_data[69][2] = 0;
        pixel_data[69][3] = 0;
        pixel_data[69][4] = 0;
        pixel_data[69][5] = 0;
        pixel_data[69][6] = 0;
        pixel_data[69][7] = 0;
        pixel_data[69][8] = 0;
        pixel_data[69][9] = 0;
        pixel_data[69][10] = 0;
        pixel_data[69][11] = 0;
        pixel_data[69][12] = 0;
        pixel_data[69][13] = 0;
        pixel_data[69][14] = 0;
        pixel_data[69][15] = 0;
        pixel_data[69][16] = 0;
        pixel_data[69][17] = 0;
        pixel_data[69][18] = 0;
        pixel_data[69][19] = 0;
        pixel_data[69][20] = 0;
        pixel_data[69][21] = 0;
        pixel_data[69][22] = 0;
        pixel_data[69][23] = 0;
        pixel_data[69][24] = 0;
        pixel_data[69][25] = 0;
        pixel_data[69][26] = 0;
        pixel_data[69][27] = 0;
        pixel_data[69][28] = 0;
        pixel_data[69][29] = 0;
        pixel_data[69][30] = 0;
        pixel_data[69][31] = 0;
        pixel_data[69][32] = 0;
        pixel_data[69][33] = 0;
        pixel_data[69][34] = 0;
        pixel_data[69][35] = 0;
        pixel_data[69][36] = 0;
        pixel_data[69][37] = 0;
        pixel_data[69][38] = 0;
        pixel_data[69][39] = 0;
        pixel_data[69][40] = 0;
        pixel_data[69][41] = 0;
        pixel_data[69][42] = 0;
        pixel_data[69][43] = 0;
        pixel_data[69][44] = 0;
        pixel_data[69][45] = 0;
        pixel_data[69][46] = 0;
        pixel_data[69][47] = 0;
        pixel_data[69][48] = 0;
        pixel_data[69][49] = 0;
        pixel_data[69][50] = 0;
        pixel_data[69][51] = 0;
        pixel_data[69][52] = 0;
        pixel_data[69][53] = 0;
        pixel_data[69][54] = 0;
        pixel_data[69][55] = 0;
        pixel_data[69][56] = 0;
        pixel_data[69][57] = 0;
        pixel_data[69][58] = 0;
        pixel_data[69][59] = 0;
        pixel_data[69][60] = 0;
        pixel_data[69][61] = 0;
        pixel_data[69][62] = 0;
        pixel_data[69][63] = 0;
        pixel_data[69][64] = 0;
        pixel_data[69][65] = 0;
        pixel_data[69][66] = 0;
        pixel_data[69][67] = 0;
        pixel_data[69][68] = 0;
        pixel_data[69][69] = 0;
        pixel_data[69][70] = 0;
        pixel_data[69][71] = 0;
        pixel_data[69][72] = 0;
        pixel_data[69][73] = 0;
        pixel_data[69][74] = 0;
        pixel_data[69][75] = 0;
        pixel_data[69][76] = 0;
        pixel_data[69][77] = 0;
        pixel_data[69][78] = 0;
        pixel_data[69][79] = 0;
        pixel_data[69][80] = 0;
        pixel_data[69][81] = 0;
        pixel_data[69][82] = 0;
        pixel_data[69][83] = 0;
        pixel_data[69][84] = 0;
        pixel_data[69][85] = 0;
        pixel_data[69][86] = 0;
        pixel_data[69][87] = 0;
        pixel_data[69][88] = 0;
        pixel_data[69][89] = 0;
        pixel_data[69][90] = 0;
        pixel_data[69][91] = 0;
        pixel_data[69][92] = 0;
        pixel_data[69][93] = 0;
        pixel_data[69][94] = 0;
        pixel_data[69][95] = 0;
        pixel_data[69][96] = 0;
        pixel_data[69][97] = 0;
        pixel_data[69][98] = 0;
        pixel_data[69][99] = 0;
        pixel_data[69][100] = 0;
        pixel_data[69][101] = 0;
        pixel_data[69][102] = 0;
        pixel_data[69][103] = 0;
        pixel_data[69][104] = 0;
        pixel_data[69][105] = 0;
        pixel_data[69][106] = 0;
        pixel_data[69][107] = 0;
        pixel_data[69][108] = 0;
        pixel_data[69][109] = 0;
        pixel_data[69][110] = 0;
        pixel_data[69][111] = 0;
        pixel_data[69][112] = 0;
        pixel_data[69][113] = 0;
        pixel_data[69][114] = 0;
        pixel_data[69][115] = 0;
        pixel_data[69][116] = 0;
        pixel_data[69][117] = 0;
        pixel_data[69][118] = 0;
        pixel_data[69][119] = 0;
        pixel_data[69][120] = 0;
        pixel_data[69][121] = 0;
        pixel_data[69][122] = 0;
        pixel_data[69][123] = 0;
        pixel_data[69][124] = 0;
        pixel_data[69][125] = 0;
        pixel_data[69][126] = 0;
        pixel_data[69][127] = 0;
        pixel_data[69][128] = 0;
        pixel_data[69][129] = 0;
        pixel_data[69][130] = 0;
        pixel_data[69][131] = 0;
        pixel_data[69][132] = 0;
        pixel_data[69][133] = 0;
        pixel_data[69][134] = 0;
        pixel_data[69][135] = 0;
        pixel_data[69][136] = 0;
        pixel_data[69][137] = 0;
        pixel_data[69][138] = 0;
        pixel_data[69][139] = 0;
        pixel_data[69][140] = 0;
        pixel_data[69][141] = 0;
        pixel_data[69][142] = 0;
        pixel_data[69][143] = 0;
        pixel_data[69][144] = 0;
        pixel_data[69][145] = 0;
        pixel_data[69][146] = 0;
        pixel_data[69][147] = 0;
        pixel_data[69][148] = 0;
        pixel_data[69][149] = 0;
        pixel_data[69][150] = 0;
        pixel_data[69][151] = 0;
        pixel_data[69][152] = 0;
        pixel_data[69][153] = 0;
        pixel_data[69][154] = 0;
        pixel_data[69][155] = 0;
        pixel_data[69][156] = 0;
        pixel_data[69][157] = 0;
        pixel_data[69][158] = 0;
        pixel_data[69][159] = 0;
        pixel_data[69][160] = 0;
        pixel_data[69][161] = 0;
        pixel_data[69][162] = 0;
        pixel_data[69][163] = 0;
        pixel_data[69][164] = 0;
        pixel_data[69][165] = 0;
        pixel_data[69][166] = 0;
        pixel_data[69][167] = 0;
        pixel_data[69][168] = 0;
        pixel_data[69][169] = 0;
        pixel_data[69][170] = 0;
        pixel_data[69][171] = 0;
        pixel_data[69][172] = 0;
        pixel_data[69][173] = 0;
        pixel_data[69][174] = 0;
        pixel_data[69][175] = 0;
        pixel_data[69][176] = 0;
        pixel_data[69][177] = 0;
        pixel_data[69][178] = 0;
        pixel_data[69][179] = 0;
        pixel_data[69][180] = 0;
        pixel_data[69][181] = 0;
        pixel_data[69][182] = 0;
        pixel_data[69][183] = 0;
        pixel_data[69][184] = 0;
        pixel_data[69][185] = 0;
        pixel_data[69][186] = 0;
        pixel_data[69][187] = 0;
        pixel_data[69][188] = 0;
        pixel_data[69][189] = 0;
        pixel_data[69][190] = 0;
        pixel_data[69][191] = 0;
        pixel_data[69][192] = 0;
        pixel_data[69][193] = 0;
        pixel_data[69][194] = 0;
        pixel_data[69][195] = 0;
        pixel_data[69][196] = 0;
        pixel_data[69][197] = 0;
        pixel_data[69][198] = 0;
        pixel_data[69][199] = 0; // y=69
        pixel_data[70][0] = 0;
        pixel_data[70][1] = 0;
        pixel_data[70][2] = 0;
        pixel_data[70][3] = 0;
        pixel_data[70][4] = 0;
        pixel_data[70][5] = 0;
        pixel_data[70][6] = 0;
        pixel_data[70][7] = 0;
        pixel_data[70][8] = 0;
        pixel_data[70][9] = 0;
        pixel_data[70][10] = 0;
        pixel_data[70][11] = 0;
        pixel_data[70][12] = 0;
        pixel_data[70][13] = 0;
        pixel_data[70][14] = 0;
        pixel_data[70][15] = 0;
        pixel_data[70][16] = 0;
        pixel_data[70][17] = 0;
        pixel_data[70][18] = 0;
        pixel_data[70][19] = 0;
        pixel_data[70][20] = 0;
        pixel_data[70][21] = 0;
        pixel_data[70][22] = 0;
        pixel_data[70][23] = 0;
        pixel_data[70][24] = 0;
        pixel_data[70][25] = 0;
        pixel_data[70][26] = 0;
        pixel_data[70][27] = 0;
        pixel_data[70][28] = 0;
        pixel_data[70][29] = 0;
        pixel_data[70][30] = 0;
        pixel_data[70][31] = 0;
        pixel_data[70][32] = 0;
        pixel_data[70][33] = 0;
        pixel_data[70][34] = 0;
        pixel_data[70][35] = 0;
        pixel_data[70][36] = 0;
        pixel_data[70][37] = 0;
        pixel_data[70][38] = 0;
        pixel_data[70][39] = 0;
        pixel_data[70][40] = 0;
        pixel_data[70][41] = 0;
        pixel_data[70][42] = 0;
        pixel_data[70][43] = 0;
        pixel_data[70][44] = 0;
        pixel_data[70][45] = 0;
        pixel_data[70][46] = 0;
        pixel_data[70][47] = 0;
        pixel_data[70][48] = 0;
        pixel_data[70][49] = 0;
        pixel_data[70][50] = 0;
        pixel_data[70][51] = 0;
        pixel_data[70][52] = 0;
        pixel_data[70][53] = 0;
        pixel_data[70][54] = 0;
        pixel_data[70][55] = 0;
        pixel_data[70][56] = 0;
        pixel_data[70][57] = 0;
        pixel_data[70][58] = 0;
        pixel_data[70][59] = 0;
        pixel_data[70][60] = 0;
        pixel_data[70][61] = 0;
        pixel_data[70][62] = 0;
        pixel_data[70][63] = 0;
        pixel_data[70][64] = 0;
        pixel_data[70][65] = 0;
        pixel_data[70][66] = 0;
        pixel_data[70][67] = 0;
        pixel_data[70][68] = 0;
        pixel_data[70][69] = 0;
        pixel_data[70][70] = 0;
        pixel_data[70][71] = 0;
        pixel_data[70][72] = 0;
        pixel_data[70][73] = 0;
        pixel_data[70][74] = 0;
        pixel_data[70][75] = 0;
        pixel_data[70][76] = 0;
        pixel_data[70][77] = 0;
        pixel_data[70][78] = 0;
        pixel_data[70][79] = 0;
        pixel_data[70][80] = 0;
        pixel_data[70][81] = 0;
        pixel_data[70][82] = 0;
        pixel_data[70][83] = 0;
        pixel_data[70][84] = 0;
        pixel_data[70][85] = 0;
        pixel_data[70][86] = 0;
        pixel_data[70][87] = 0;
        pixel_data[70][88] = 0;
        pixel_data[70][89] = 0;
        pixel_data[70][90] = 0;
        pixel_data[70][91] = 0;
        pixel_data[70][92] = 0;
        pixel_data[70][93] = 0;
        pixel_data[70][94] = 0;
        pixel_data[70][95] = 0;
        pixel_data[70][96] = 0;
        pixel_data[70][97] = 0;
        pixel_data[70][98] = 0;
        pixel_data[70][99] = 0;
        pixel_data[70][100] = 0;
        pixel_data[70][101] = 0;
        pixel_data[70][102] = 0;
        pixel_data[70][103] = 0;
        pixel_data[70][104] = 0;
        pixel_data[70][105] = 0;
        pixel_data[70][106] = 0;
        pixel_data[70][107] = 0;
        pixel_data[70][108] = 0;
        pixel_data[70][109] = 0;
        pixel_data[70][110] = 0;
        pixel_data[70][111] = 0;
        pixel_data[70][112] = 0;
        pixel_data[70][113] = 0;
        pixel_data[70][114] = 0;
        pixel_data[70][115] = 0;
        pixel_data[70][116] = 0;
        pixel_data[70][117] = 0;
        pixel_data[70][118] = 0;
        pixel_data[70][119] = 0;
        pixel_data[70][120] = 0;
        pixel_data[70][121] = 0;
        pixel_data[70][122] = 0;
        pixel_data[70][123] = 0;
        pixel_data[70][124] = 0;
        pixel_data[70][125] = 0;
        pixel_data[70][126] = 0;
        pixel_data[70][127] = 0;
        pixel_data[70][128] = 0;
        pixel_data[70][129] = 0;
        pixel_data[70][130] = 0;
        pixel_data[70][131] = 0;
        pixel_data[70][132] = 0;
        pixel_data[70][133] = 0;
        pixel_data[70][134] = 0;
        pixel_data[70][135] = 0;
        pixel_data[70][136] = 0;
        pixel_data[70][137] = 0;
        pixel_data[70][138] = 0;
        pixel_data[70][139] = 0;
        pixel_data[70][140] = 0;
        pixel_data[70][141] = 0;
        pixel_data[70][142] = 0;
        pixel_data[70][143] = 0;
        pixel_data[70][144] = 0;
        pixel_data[70][145] = 0;
        pixel_data[70][146] = 0;
        pixel_data[70][147] = 0;
        pixel_data[70][148] = 0;
        pixel_data[70][149] = 0;
        pixel_data[70][150] = 0;
        pixel_data[70][151] = 0;
        pixel_data[70][152] = 0;
        pixel_data[70][153] = 0;
        pixel_data[70][154] = 0;
        pixel_data[70][155] = 0;
        pixel_data[70][156] = 0;
        pixel_data[70][157] = 0;
        pixel_data[70][158] = 0;
        pixel_data[70][159] = 0;
        pixel_data[70][160] = 0;
        pixel_data[70][161] = 0;
        pixel_data[70][162] = 0;
        pixel_data[70][163] = 0;
        pixel_data[70][164] = 0;
        pixel_data[70][165] = 0;
        pixel_data[70][166] = 0;
        pixel_data[70][167] = 0;
        pixel_data[70][168] = 0;
        pixel_data[70][169] = 0;
        pixel_data[70][170] = 0;
        pixel_data[70][171] = 0;
        pixel_data[70][172] = 0;
        pixel_data[70][173] = 0;
        pixel_data[70][174] = 0;
        pixel_data[70][175] = 0;
        pixel_data[70][176] = 0;
        pixel_data[70][177] = 0;
        pixel_data[70][178] = 0;
        pixel_data[70][179] = 0;
        pixel_data[70][180] = 0;
        pixel_data[70][181] = 0;
        pixel_data[70][182] = 0;
        pixel_data[70][183] = 0;
        pixel_data[70][184] = 0;
        pixel_data[70][185] = 0;
        pixel_data[70][186] = 0;
        pixel_data[70][187] = 0;
        pixel_data[70][188] = 0;
        pixel_data[70][189] = 0;
        pixel_data[70][190] = 0;
        pixel_data[70][191] = 0;
        pixel_data[70][192] = 0;
        pixel_data[70][193] = 0;
        pixel_data[70][194] = 0;
        pixel_data[70][195] = 0;
        pixel_data[70][196] = 0;
        pixel_data[70][197] = 0;
        pixel_data[70][198] = 0;
        pixel_data[70][199] = 0; // y=70
        pixel_data[71][0] = 0;
        pixel_data[71][1] = 0;
        pixel_data[71][2] = 0;
        pixel_data[71][3] = 0;
        pixel_data[71][4] = 0;
        pixel_data[71][5] = 0;
        pixel_data[71][6] = 0;
        pixel_data[71][7] = 0;
        pixel_data[71][8] = 0;
        pixel_data[71][9] = 0;
        pixel_data[71][10] = 0;
        pixel_data[71][11] = 0;
        pixel_data[71][12] = 0;
        pixel_data[71][13] = 0;
        pixel_data[71][14] = 0;
        pixel_data[71][15] = 0;
        pixel_data[71][16] = 0;
        pixel_data[71][17] = 0;
        pixel_data[71][18] = 0;
        pixel_data[71][19] = 0;
        pixel_data[71][20] = 0;
        pixel_data[71][21] = 0;
        pixel_data[71][22] = 0;
        pixel_data[71][23] = 0;
        pixel_data[71][24] = 0;
        pixel_data[71][25] = 0;
        pixel_data[71][26] = 0;
        pixel_data[71][27] = 0;
        pixel_data[71][28] = 0;
        pixel_data[71][29] = 0;
        pixel_data[71][30] = 0;
        pixel_data[71][31] = 0;
        pixel_data[71][32] = 0;
        pixel_data[71][33] = 0;
        pixel_data[71][34] = 0;
        pixel_data[71][35] = 0;
        pixel_data[71][36] = 0;
        pixel_data[71][37] = 0;
        pixel_data[71][38] = 0;
        pixel_data[71][39] = 0;
        pixel_data[71][40] = 0;
        pixel_data[71][41] = 0;
        pixel_data[71][42] = 0;
        pixel_data[71][43] = 0;
        pixel_data[71][44] = 0;
        pixel_data[71][45] = 0;
        pixel_data[71][46] = 0;
        pixel_data[71][47] = 0;
        pixel_data[71][48] = 0;
        pixel_data[71][49] = 0;
        pixel_data[71][50] = 0;
        pixel_data[71][51] = 0;
        pixel_data[71][52] = 0;
        pixel_data[71][53] = 0;
        pixel_data[71][54] = 0;
        pixel_data[71][55] = 0;
        pixel_data[71][56] = 0;
        pixel_data[71][57] = 0;
        pixel_data[71][58] = 0;
        pixel_data[71][59] = 0;
        pixel_data[71][60] = 0;
        pixel_data[71][61] = 0;
        pixel_data[71][62] = 0;
        pixel_data[71][63] = 0;
        pixel_data[71][64] = 0;
        pixel_data[71][65] = 0;
        pixel_data[71][66] = 0;
        pixel_data[71][67] = 0;
        pixel_data[71][68] = 0;
        pixel_data[71][69] = 0;
        pixel_data[71][70] = 0;
        pixel_data[71][71] = 0;
        pixel_data[71][72] = 0;
        pixel_data[71][73] = 0;
        pixel_data[71][74] = 0;
        pixel_data[71][75] = 0;
        pixel_data[71][76] = 0;
        pixel_data[71][77] = 0;
        pixel_data[71][78] = 0;
        pixel_data[71][79] = 0;
        pixel_data[71][80] = 0;
        pixel_data[71][81] = 0;
        pixel_data[71][82] = 0;
        pixel_data[71][83] = 0;
        pixel_data[71][84] = 0;
        pixel_data[71][85] = 0;
        pixel_data[71][86] = 0;
        pixel_data[71][87] = 0;
        pixel_data[71][88] = 0;
        pixel_data[71][89] = 0;
        pixel_data[71][90] = 0;
        pixel_data[71][91] = 0;
        pixel_data[71][92] = 0;
        pixel_data[71][93] = 0;
        pixel_data[71][94] = 0;
        pixel_data[71][95] = 0;
        pixel_data[71][96] = 0;
        pixel_data[71][97] = 0;
        pixel_data[71][98] = 0;
        pixel_data[71][99] = 0;
        pixel_data[71][100] = 0;
        pixel_data[71][101] = 0;
        pixel_data[71][102] = 0;
        pixel_data[71][103] = 0;
        pixel_data[71][104] = 0;
        pixel_data[71][105] = 0;
        pixel_data[71][106] = 0;
        pixel_data[71][107] = 0;
        pixel_data[71][108] = 0;
        pixel_data[71][109] = 0;
        pixel_data[71][110] = 0;
        pixel_data[71][111] = 0;
        pixel_data[71][112] = 0;
        pixel_data[71][113] = 0;
        pixel_data[71][114] = 0;
        pixel_data[71][115] = 0;
        pixel_data[71][116] = 0;
        pixel_data[71][117] = 0;
        pixel_data[71][118] = 0;
        pixel_data[71][119] = 0;
        pixel_data[71][120] = 0;
        pixel_data[71][121] = 0;
        pixel_data[71][122] = 0;
        pixel_data[71][123] = 0;
        pixel_data[71][124] = 0;
        pixel_data[71][125] = 0;
        pixel_data[71][126] = 0;
        pixel_data[71][127] = 0;
        pixel_data[71][128] = 0;
        pixel_data[71][129] = 0;
        pixel_data[71][130] = 0;
        pixel_data[71][131] = 0;
        pixel_data[71][132] = 0;
        pixel_data[71][133] = 0;
        pixel_data[71][134] = 0;
        pixel_data[71][135] = 0;
        pixel_data[71][136] = 0;
        pixel_data[71][137] = 0;
        pixel_data[71][138] = 0;
        pixel_data[71][139] = 0;
        pixel_data[71][140] = 0;
        pixel_data[71][141] = 0;
        pixel_data[71][142] = 0;
        pixel_data[71][143] = 0;
        pixel_data[71][144] = 0;
        pixel_data[71][145] = 0;
        pixel_data[71][146] = 0;
        pixel_data[71][147] = 0;
        pixel_data[71][148] = 0;
        pixel_data[71][149] = 0;
        pixel_data[71][150] = 0;
        pixel_data[71][151] = 0;
        pixel_data[71][152] = 0;
        pixel_data[71][153] = 0;
        pixel_data[71][154] = 0;
        pixel_data[71][155] = 0;
        pixel_data[71][156] = 0;
        pixel_data[71][157] = 0;
        pixel_data[71][158] = 0;
        pixel_data[71][159] = 0;
        pixel_data[71][160] = 0;
        pixel_data[71][161] = 0;
        pixel_data[71][162] = 0;
        pixel_data[71][163] = 0;
        pixel_data[71][164] = 0;
        pixel_data[71][165] = 0;
        pixel_data[71][166] = 0;
        pixel_data[71][167] = 0;
        pixel_data[71][168] = 0;
        pixel_data[71][169] = 0;
        pixel_data[71][170] = 0;
        pixel_data[71][171] = 0;
        pixel_data[71][172] = 0;
        pixel_data[71][173] = 0;
        pixel_data[71][174] = 0;
        pixel_data[71][175] = 0;
        pixel_data[71][176] = 0;
        pixel_data[71][177] = 0;
        pixel_data[71][178] = 0;
        pixel_data[71][179] = 0;
        pixel_data[71][180] = 0;
        pixel_data[71][181] = 0;
        pixel_data[71][182] = 0;
        pixel_data[71][183] = 0;
        pixel_data[71][184] = 0;
        pixel_data[71][185] = 0;
        pixel_data[71][186] = 0;
        pixel_data[71][187] = 0;
        pixel_data[71][188] = 0;
        pixel_data[71][189] = 0;
        pixel_data[71][190] = 0;
        pixel_data[71][191] = 0;
        pixel_data[71][192] = 0;
        pixel_data[71][193] = 0;
        pixel_data[71][194] = 0;
        pixel_data[71][195] = 0;
        pixel_data[71][196] = 0;
        pixel_data[71][197] = 0;
        pixel_data[71][198] = 0;
        pixel_data[71][199] = 0; // y=71
        pixel_data[72][0] = 0;
        pixel_data[72][1] = 0;
        pixel_data[72][2] = 0;
        pixel_data[72][3] = 0;
        pixel_data[72][4] = 0;
        pixel_data[72][5] = 0;
        pixel_data[72][6] = 0;
        pixel_data[72][7] = 0;
        pixel_data[72][8] = 0;
        pixel_data[72][9] = 0;
        pixel_data[72][10] = 0;
        pixel_data[72][11] = 0;
        pixel_data[72][12] = 0;
        pixel_data[72][13] = 0;
        pixel_data[72][14] = 0;
        pixel_data[72][15] = 0;
        pixel_data[72][16] = 0;
        pixel_data[72][17] = 0;
        pixel_data[72][18] = 0;
        pixel_data[72][19] = 0;
        pixel_data[72][20] = 0;
        pixel_data[72][21] = 0;
        pixel_data[72][22] = 0;
        pixel_data[72][23] = 0;
        pixel_data[72][24] = 0;
        pixel_data[72][25] = 0;
        pixel_data[72][26] = 0;
        pixel_data[72][27] = 0;
        pixel_data[72][28] = 0;
        pixel_data[72][29] = 0;
        pixel_data[72][30] = 0;
        pixel_data[72][31] = 0;
        pixel_data[72][32] = 0;
        pixel_data[72][33] = 0;
        pixel_data[72][34] = 0;
        pixel_data[72][35] = 0;
        pixel_data[72][36] = 0;
        pixel_data[72][37] = 0;
        pixel_data[72][38] = 0;
        pixel_data[72][39] = 0;
        pixel_data[72][40] = 0;
        pixel_data[72][41] = 0;
        pixel_data[72][42] = 0;
        pixel_data[72][43] = 0;
        pixel_data[72][44] = 0;
        pixel_data[72][45] = 0;
        pixel_data[72][46] = 0;
        pixel_data[72][47] = 0;
        pixel_data[72][48] = 0;
        pixel_data[72][49] = 0;
        pixel_data[72][50] = 0;
        pixel_data[72][51] = 0;
        pixel_data[72][52] = 0;
        pixel_data[72][53] = 0;
        pixel_data[72][54] = 0;
        pixel_data[72][55] = 0;
        pixel_data[72][56] = 0;
        pixel_data[72][57] = 0;
        pixel_data[72][58] = 0;
        pixel_data[72][59] = 0;
        pixel_data[72][60] = 0;
        pixel_data[72][61] = 0;
        pixel_data[72][62] = 0;
        pixel_data[72][63] = 0;
        pixel_data[72][64] = 0;
        pixel_data[72][65] = 0;
        pixel_data[72][66] = 0;
        pixel_data[72][67] = 0;
        pixel_data[72][68] = 0;
        pixel_data[72][69] = 0;
        pixel_data[72][70] = 0;
        pixel_data[72][71] = 0;
        pixel_data[72][72] = 0;
        pixel_data[72][73] = 0;
        pixel_data[72][74] = 0;
        pixel_data[72][75] = 0;
        pixel_data[72][76] = 0;
        pixel_data[72][77] = 0;
        pixel_data[72][78] = 0;
        pixel_data[72][79] = 0;
        pixel_data[72][80] = 0;
        pixel_data[72][81] = 0;
        pixel_data[72][82] = 0;
        pixel_data[72][83] = 0;
        pixel_data[72][84] = 0;
        pixel_data[72][85] = 0;
        pixel_data[72][86] = 0;
        pixel_data[72][87] = 0;
        pixel_data[72][88] = 0;
        pixel_data[72][89] = 0;
        pixel_data[72][90] = 0;
        pixel_data[72][91] = 0;
        pixel_data[72][92] = 0;
        pixel_data[72][93] = 0;
        pixel_data[72][94] = 0;
        pixel_data[72][95] = 0;
        pixel_data[72][96] = 0;
        pixel_data[72][97] = 0;
        pixel_data[72][98] = 0;
        pixel_data[72][99] = 0;
        pixel_data[72][100] = 0;
        pixel_data[72][101] = 0;
        pixel_data[72][102] = 0;
        pixel_data[72][103] = 0;
        pixel_data[72][104] = 0;
        pixel_data[72][105] = 0;
        pixel_data[72][106] = 0;
        pixel_data[72][107] = 0;
        pixel_data[72][108] = 0;
        pixel_data[72][109] = 0;
        pixel_data[72][110] = 0;
        pixel_data[72][111] = 0;
        pixel_data[72][112] = 0;
        pixel_data[72][113] = 0;
        pixel_data[72][114] = 0;
        pixel_data[72][115] = 0;
        pixel_data[72][116] = 0;
        pixel_data[72][117] = 0;
        pixel_data[72][118] = 0;
        pixel_data[72][119] = 0;
        pixel_data[72][120] = 0;
        pixel_data[72][121] = 0;
        pixel_data[72][122] = 0;
        pixel_data[72][123] = 0;
        pixel_data[72][124] = 0;
        pixel_data[72][125] = 0;
        pixel_data[72][126] = 0;
        pixel_data[72][127] = 0;
        pixel_data[72][128] = 0;
        pixel_data[72][129] = 0;
        pixel_data[72][130] = 0;
        pixel_data[72][131] = 0;
        pixel_data[72][132] = 0;
        pixel_data[72][133] = 0;
        pixel_data[72][134] = 0;
        pixel_data[72][135] = 0;
        pixel_data[72][136] = 0;
        pixel_data[72][137] = 0;
        pixel_data[72][138] = 0;
        pixel_data[72][139] = 0;
        pixel_data[72][140] = 0;
        pixel_data[72][141] = 0;
        pixel_data[72][142] = 0;
        pixel_data[72][143] = 0;
        pixel_data[72][144] = 0;
        pixel_data[72][145] = 0;
        pixel_data[72][146] = 0;
        pixel_data[72][147] = 0;
        pixel_data[72][148] = 0;
        pixel_data[72][149] = 0;
        pixel_data[72][150] = 0;
        pixel_data[72][151] = 0;
        pixel_data[72][152] = 0;
        pixel_data[72][153] = 0;
        pixel_data[72][154] = 0;
        pixel_data[72][155] = 0;
        pixel_data[72][156] = 0;
        pixel_data[72][157] = 0;
        pixel_data[72][158] = 0;
        pixel_data[72][159] = 0;
        pixel_data[72][160] = 0;
        pixel_data[72][161] = 0;
        pixel_data[72][162] = 0;
        pixel_data[72][163] = 0;
        pixel_data[72][164] = 0;
        pixel_data[72][165] = 0;
        pixel_data[72][166] = 0;
        pixel_data[72][167] = 0;
        pixel_data[72][168] = 0;
        pixel_data[72][169] = 0;
        pixel_data[72][170] = 0;
        pixel_data[72][171] = 0;
        pixel_data[72][172] = 0;
        pixel_data[72][173] = 0;
        pixel_data[72][174] = 0;
        pixel_data[72][175] = 0;
        pixel_data[72][176] = 0;
        pixel_data[72][177] = 0;
        pixel_data[72][178] = 0;
        pixel_data[72][179] = 0;
        pixel_data[72][180] = 0;
        pixel_data[72][181] = 0;
        pixel_data[72][182] = 0;
        pixel_data[72][183] = 0;
        pixel_data[72][184] = 0;
        pixel_data[72][185] = 0;
        pixel_data[72][186] = 0;
        pixel_data[72][187] = 0;
        pixel_data[72][188] = 0;
        pixel_data[72][189] = 0;
        pixel_data[72][190] = 0;
        pixel_data[72][191] = 0;
        pixel_data[72][192] = 0;
        pixel_data[72][193] = 0;
        pixel_data[72][194] = 0;
        pixel_data[72][195] = 0;
        pixel_data[72][196] = 0;
        pixel_data[72][197] = 0;
        pixel_data[72][198] = 0;
        pixel_data[72][199] = 0; // y=72
        pixel_data[73][0] = 0;
        pixel_data[73][1] = 0;
        pixel_data[73][2] = 0;
        pixel_data[73][3] = 0;
        pixel_data[73][4] = 0;
        pixel_data[73][5] = 0;
        pixel_data[73][6] = 0;
        pixel_data[73][7] = 0;
        pixel_data[73][8] = 0;
        pixel_data[73][9] = 0;
        pixel_data[73][10] = 0;
        pixel_data[73][11] = 0;
        pixel_data[73][12] = 0;
        pixel_data[73][13] = 0;
        pixel_data[73][14] = 0;
        pixel_data[73][15] = 0;
        pixel_data[73][16] = 0;
        pixel_data[73][17] = 0;
        pixel_data[73][18] = 0;
        pixel_data[73][19] = 0;
        pixel_data[73][20] = 0;
        pixel_data[73][21] = 0;
        pixel_data[73][22] = 0;
        pixel_data[73][23] = 0;
        pixel_data[73][24] = 0;
        pixel_data[73][25] = 0;
        pixel_data[73][26] = 0;
        pixel_data[73][27] = 0;
        pixel_data[73][28] = 0;
        pixel_data[73][29] = 0;
        pixel_data[73][30] = 0;
        pixel_data[73][31] = 0;
        pixel_data[73][32] = 0;
        pixel_data[73][33] = 0;
        pixel_data[73][34] = 0;
        pixel_data[73][35] = 0;
        pixel_data[73][36] = 0;
        pixel_data[73][37] = 0;
        pixel_data[73][38] = 0;
        pixel_data[73][39] = 0;
        pixel_data[73][40] = 0;
        pixel_data[73][41] = 0;
        pixel_data[73][42] = 0;
        pixel_data[73][43] = 0;
        pixel_data[73][44] = 0;
        pixel_data[73][45] = 0;
        pixel_data[73][46] = 0;
        pixel_data[73][47] = 0;
        pixel_data[73][48] = 0;
        pixel_data[73][49] = 0;
        pixel_data[73][50] = 0;
        pixel_data[73][51] = 0;
        pixel_data[73][52] = 0;
        pixel_data[73][53] = 0;
        pixel_data[73][54] = 0;
        pixel_data[73][55] = 0;
        pixel_data[73][56] = 0;
        pixel_data[73][57] = 0;
        pixel_data[73][58] = 0;
        pixel_data[73][59] = 0;
        pixel_data[73][60] = 0;
        pixel_data[73][61] = 0;
        pixel_data[73][62] = 0;
        pixel_data[73][63] = 0;
        pixel_data[73][64] = 0;
        pixel_data[73][65] = 0;
        pixel_data[73][66] = 0;
        pixel_data[73][67] = 0;
        pixel_data[73][68] = 0;
        pixel_data[73][69] = 0;
        pixel_data[73][70] = 0;
        pixel_data[73][71] = 0;
        pixel_data[73][72] = 0;
        pixel_data[73][73] = 0;
        pixel_data[73][74] = 0;
        pixel_data[73][75] = 0;
        pixel_data[73][76] = 0;
        pixel_data[73][77] = 0;
        pixel_data[73][78] = 0;
        pixel_data[73][79] = 0;
        pixel_data[73][80] = 0;
        pixel_data[73][81] = 0;
        pixel_data[73][82] = 0;
        pixel_data[73][83] = 0;
        pixel_data[73][84] = 0;
        pixel_data[73][85] = 0;
        pixel_data[73][86] = 0;
        pixel_data[73][87] = 0;
        pixel_data[73][88] = 0;
        pixel_data[73][89] = 0;
        pixel_data[73][90] = 0;
        pixel_data[73][91] = 0;
        pixel_data[73][92] = 0;
        pixel_data[73][93] = 0;
        pixel_data[73][94] = 0;
        pixel_data[73][95] = 0;
        pixel_data[73][96] = 0;
        pixel_data[73][97] = 0;
        pixel_data[73][98] = 0;
        pixel_data[73][99] = 0;
        pixel_data[73][100] = 0;
        pixel_data[73][101] = 0;
        pixel_data[73][102] = 0;
        pixel_data[73][103] = 0;
        pixel_data[73][104] = 0;
        pixel_data[73][105] = 0;
        pixel_data[73][106] = 0;
        pixel_data[73][107] = 0;
        pixel_data[73][108] = 0;
        pixel_data[73][109] = 0;
        pixel_data[73][110] = 0;
        pixel_data[73][111] = 0;
        pixel_data[73][112] = 0;
        pixel_data[73][113] = 0;
        pixel_data[73][114] = 0;
        pixel_data[73][115] = 0;
        pixel_data[73][116] = 0;
        pixel_data[73][117] = 0;
        pixel_data[73][118] = 0;
        pixel_data[73][119] = 0;
        pixel_data[73][120] = 0;
        pixel_data[73][121] = 0;
        pixel_data[73][122] = 0;
        pixel_data[73][123] = 0;
        pixel_data[73][124] = 0;
        pixel_data[73][125] = 0;
        pixel_data[73][126] = 0;
        pixel_data[73][127] = 0;
        pixel_data[73][128] = 0;
        pixel_data[73][129] = 0;
        pixel_data[73][130] = 0;
        pixel_data[73][131] = 0;
        pixel_data[73][132] = 0;
        pixel_data[73][133] = 0;
        pixel_data[73][134] = 0;
        pixel_data[73][135] = 0;
        pixel_data[73][136] = 0;
        pixel_data[73][137] = 0;
        pixel_data[73][138] = 0;
        pixel_data[73][139] = 0;
        pixel_data[73][140] = 0;
        pixel_data[73][141] = 0;
        pixel_data[73][142] = 0;
        pixel_data[73][143] = 0;
        pixel_data[73][144] = 0;
        pixel_data[73][145] = 0;
        pixel_data[73][146] = 0;
        pixel_data[73][147] = 0;
        pixel_data[73][148] = 0;
        pixel_data[73][149] = 0;
        pixel_data[73][150] = 0;
        pixel_data[73][151] = 0;
        pixel_data[73][152] = 0;
        pixel_data[73][153] = 0;
        pixel_data[73][154] = 0;
        pixel_data[73][155] = 0;
        pixel_data[73][156] = 0;
        pixel_data[73][157] = 0;
        pixel_data[73][158] = 0;
        pixel_data[73][159] = 0;
        pixel_data[73][160] = 0;
        pixel_data[73][161] = 0;
        pixel_data[73][162] = 0;
        pixel_data[73][163] = 0;
        pixel_data[73][164] = 0;
        pixel_data[73][165] = 0;
        pixel_data[73][166] = 0;
        pixel_data[73][167] = 0;
        pixel_data[73][168] = 0;
        pixel_data[73][169] = 0;
        pixel_data[73][170] = 0;
        pixel_data[73][171] = 0;
        pixel_data[73][172] = 0;
        pixel_data[73][173] = 0;
        pixel_data[73][174] = 0;
        pixel_data[73][175] = 0;
        pixel_data[73][176] = 0;
        pixel_data[73][177] = 0;
        pixel_data[73][178] = 0;
        pixel_data[73][179] = 0;
        pixel_data[73][180] = 0;
        pixel_data[73][181] = 0;
        pixel_data[73][182] = 0;
        pixel_data[73][183] = 0;
        pixel_data[73][184] = 0;
        pixel_data[73][185] = 0;
        pixel_data[73][186] = 0;
        pixel_data[73][187] = 0;
        pixel_data[73][188] = 0;
        pixel_data[73][189] = 0;
        pixel_data[73][190] = 0;
        pixel_data[73][191] = 0;
        pixel_data[73][192] = 0;
        pixel_data[73][193] = 0;
        pixel_data[73][194] = 0;
        pixel_data[73][195] = 0;
        pixel_data[73][196] = 0;
        pixel_data[73][197] = 0;
        pixel_data[73][198] = 0;
        pixel_data[73][199] = 0; // y=73
        pixel_data[74][0] = 0;
        pixel_data[74][1] = 0;
        pixel_data[74][2] = 0;
        pixel_data[74][3] = 0;
        pixel_data[74][4] = 0;
        pixel_data[74][5] = 0;
        pixel_data[74][6] = 0;
        pixel_data[74][7] = 0;
        pixel_data[74][8] = 0;
        pixel_data[74][9] = 0;
        pixel_data[74][10] = 0;
        pixel_data[74][11] = 0;
        pixel_data[74][12] = 0;
        pixel_data[74][13] = 0;
        pixel_data[74][14] = 0;
        pixel_data[74][15] = 0;
        pixel_data[74][16] = 0;
        pixel_data[74][17] = 0;
        pixel_data[74][18] = 0;
        pixel_data[74][19] = 0;
        pixel_data[74][20] = 0;
        pixel_data[74][21] = 0;
        pixel_data[74][22] = 0;
        pixel_data[74][23] = 0;
        pixel_data[74][24] = 0;
        pixel_data[74][25] = 0;
        pixel_data[74][26] = 0;
        pixel_data[74][27] = 0;
        pixel_data[74][28] = 0;
        pixel_data[74][29] = 0;
        pixel_data[74][30] = 0;
        pixel_data[74][31] = 0;
        pixel_data[74][32] = 0;
        pixel_data[74][33] = 0;
        pixel_data[74][34] = 0;
        pixel_data[74][35] = 0;
        pixel_data[74][36] = 0;
        pixel_data[74][37] = 0;
        pixel_data[74][38] = 0;
        pixel_data[74][39] = 0;
        pixel_data[74][40] = 0;
        pixel_data[74][41] = 0;
        pixel_data[74][42] = 0;
        pixel_data[74][43] = 0;
        pixel_data[74][44] = 0;
        pixel_data[74][45] = 0;
        pixel_data[74][46] = 0;
        pixel_data[74][47] = 0;
        pixel_data[74][48] = 0;
        pixel_data[74][49] = 0;
        pixel_data[74][50] = 0;
        pixel_data[74][51] = 0;
        pixel_data[74][52] = 0;
        pixel_data[74][53] = 0;
        pixel_data[74][54] = 0;
        pixel_data[74][55] = 0;
        pixel_data[74][56] = 0;
        pixel_data[74][57] = 0;
        pixel_data[74][58] = 0;
        pixel_data[74][59] = 0;
        pixel_data[74][60] = 0;
        pixel_data[74][61] = 0;
        pixel_data[74][62] = 0;
        pixel_data[74][63] = 0;
        pixel_data[74][64] = 0;
        pixel_data[74][65] = 0;
        pixel_data[74][66] = 0;
        pixel_data[74][67] = 0;
        pixel_data[74][68] = 0;
        pixel_data[74][69] = 0;
        pixel_data[74][70] = 0;
        pixel_data[74][71] = 0;
        pixel_data[74][72] = 0;
        pixel_data[74][73] = 0;
        pixel_data[74][74] = 0;
        pixel_data[74][75] = 0;
        pixel_data[74][76] = 0;
        pixel_data[74][77] = 0;
        pixel_data[74][78] = 0;
        pixel_data[74][79] = 0;
        pixel_data[74][80] = 0;
        pixel_data[74][81] = 0;
        pixel_data[74][82] = 0;
        pixel_data[74][83] = 0;
        pixel_data[74][84] = 0;
        pixel_data[74][85] = 0;
        pixel_data[74][86] = 0;
        pixel_data[74][87] = 0;
        pixel_data[74][88] = 0;
        pixel_data[74][89] = 0;
        pixel_data[74][90] = 0;
        pixel_data[74][91] = 0;
        pixel_data[74][92] = 0;
        pixel_data[74][93] = 0;
        pixel_data[74][94] = 0;
        pixel_data[74][95] = 0;
        pixel_data[74][96] = 0;
        pixel_data[74][97] = 0;
        pixel_data[74][98] = 0;
        pixel_data[74][99] = 0;
        pixel_data[74][100] = 0;
        pixel_data[74][101] = 0;
        pixel_data[74][102] = 0;
        pixel_data[74][103] = 0;
        pixel_data[74][104] = 0;
        pixel_data[74][105] = 0;
        pixel_data[74][106] = 0;
        pixel_data[74][107] = 0;
        pixel_data[74][108] = 0;
        pixel_data[74][109] = 0;
        pixel_data[74][110] = 0;
        pixel_data[74][111] = 0;
        pixel_data[74][112] = 0;
        pixel_data[74][113] = 0;
        pixel_data[74][114] = 0;
        pixel_data[74][115] = 0;
        pixel_data[74][116] = 0;
        pixel_data[74][117] = 0;
        pixel_data[74][118] = 0;
        pixel_data[74][119] = 0;
        pixel_data[74][120] = 0;
        pixel_data[74][121] = 0;
        pixel_data[74][122] = 0;
        pixel_data[74][123] = 0;
        pixel_data[74][124] = 0;
        pixel_data[74][125] = 0;
        pixel_data[74][126] = 0;
        pixel_data[74][127] = 0;
        pixel_data[74][128] = 0;
        pixel_data[74][129] = 0;
        pixel_data[74][130] = 0;
        pixel_data[74][131] = 0;
        pixel_data[74][132] = 0;
        pixel_data[74][133] = 0;
        pixel_data[74][134] = 0;
        pixel_data[74][135] = 0;
        pixel_data[74][136] = 0;
        pixel_data[74][137] = 0;
        pixel_data[74][138] = 0;
        pixel_data[74][139] = 0;
        pixel_data[74][140] = 0;
        pixel_data[74][141] = 0;
        pixel_data[74][142] = 0;
        pixel_data[74][143] = 0;
        pixel_data[74][144] = 0;
        pixel_data[74][145] = 0;
        pixel_data[74][146] = 0;
        pixel_data[74][147] = 0;
        pixel_data[74][148] = 0;
        pixel_data[74][149] = 0;
        pixel_data[74][150] = 0;
        pixel_data[74][151] = 0;
        pixel_data[74][152] = 0;
        pixel_data[74][153] = 0;
        pixel_data[74][154] = 0;
        pixel_data[74][155] = 0;
        pixel_data[74][156] = 0;
        pixel_data[74][157] = 0;
        pixel_data[74][158] = 0;
        pixel_data[74][159] = 0;
        pixel_data[74][160] = 0;
        pixel_data[74][161] = 0;
        pixel_data[74][162] = 0;
        pixel_data[74][163] = 0;
        pixel_data[74][164] = 0;
        pixel_data[74][165] = 0;
        pixel_data[74][166] = 0;
        pixel_data[74][167] = 0;
        pixel_data[74][168] = 0;
        pixel_data[74][169] = 0;
        pixel_data[74][170] = 0;
        pixel_data[74][171] = 0;
        pixel_data[74][172] = 0;
        pixel_data[74][173] = 0;
        pixel_data[74][174] = 0;
        pixel_data[74][175] = 0;
        pixel_data[74][176] = 0;
        pixel_data[74][177] = 0;
        pixel_data[74][178] = 0;
        pixel_data[74][179] = 0;
        pixel_data[74][180] = 0;
        pixel_data[74][181] = 0;
        pixel_data[74][182] = 0;
        pixel_data[74][183] = 0;
        pixel_data[74][184] = 0;
        pixel_data[74][185] = 0;
        pixel_data[74][186] = 0;
        pixel_data[74][187] = 0;
        pixel_data[74][188] = 0;
        pixel_data[74][189] = 0;
        pixel_data[74][190] = 0;
        pixel_data[74][191] = 0;
        pixel_data[74][192] = 0;
        pixel_data[74][193] = 0;
        pixel_data[74][194] = 0;
        pixel_data[74][195] = 0;
        pixel_data[74][196] = 0;
        pixel_data[74][197] = 0;
        pixel_data[74][198] = 0;
        pixel_data[74][199] = 0; // y=74
        pixel_data[75][0] = 0;
        pixel_data[75][1] = 0;
        pixel_data[75][2] = 0;
        pixel_data[75][3] = 0;
        pixel_data[75][4] = 0;
        pixel_data[75][5] = 0;
        pixel_data[75][6] = 0;
        pixel_data[75][7] = 0;
        pixel_data[75][8] = 0;
        pixel_data[75][9] = 0;
        pixel_data[75][10] = 0;
        pixel_data[75][11] = 0;
        pixel_data[75][12] = 0;
        pixel_data[75][13] = 0;
        pixel_data[75][14] = 0;
        pixel_data[75][15] = 0;
        pixel_data[75][16] = 0;
        pixel_data[75][17] = 0;
        pixel_data[75][18] = 0;
        pixel_data[75][19] = 0;
        pixel_data[75][20] = 0;
        pixel_data[75][21] = 0;
        pixel_data[75][22] = 0;
        pixel_data[75][23] = 0;
        pixel_data[75][24] = 0;
        pixel_data[75][25] = 0;
        pixel_data[75][26] = 0;
        pixel_data[75][27] = 0;
        pixel_data[75][28] = 0;
        pixel_data[75][29] = 0;
        pixel_data[75][30] = 0;
        pixel_data[75][31] = 0;
        pixel_data[75][32] = 0;
        pixel_data[75][33] = 0;
        pixel_data[75][34] = 0;
        pixel_data[75][35] = 0;
        pixel_data[75][36] = 0;
        pixel_data[75][37] = 0;
        pixel_data[75][38] = 0;
        pixel_data[75][39] = 0;
        pixel_data[75][40] = 0;
        pixel_data[75][41] = 0;
        pixel_data[75][42] = 0;
        pixel_data[75][43] = 0;
        pixel_data[75][44] = 0;
        pixel_data[75][45] = 0;
        pixel_data[75][46] = 0;
        pixel_data[75][47] = 0;
        pixel_data[75][48] = 0;
        pixel_data[75][49] = 0;
        pixel_data[75][50] = 0;
        pixel_data[75][51] = 0;
        pixel_data[75][52] = 0;
        pixel_data[75][53] = 0;
        pixel_data[75][54] = 0;
        pixel_data[75][55] = 0;
        pixel_data[75][56] = 0;
        pixel_data[75][57] = 0;
        pixel_data[75][58] = 0;
        pixel_data[75][59] = 0;
        pixel_data[75][60] = 0;
        pixel_data[75][61] = 0;
        pixel_data[75][62] = 0;
        pixel_data[75][63] = 0;
        pixel_data[75][64] = 0;
        pixel_data[75][65] = 0;
        pixel_data[75][66] = 0;
        pixel_data[75][67] = 0;
        pixel_data[75][68] = 0;
        pixel_data[75][69] = 0;
        pixel_data[75][70] = 0;
        pixel_data[75][71] = 0;
        pixel_data[75][72] = 0;
        pixel_data[75][73] = 0;
        pixel_data[75][74] = 0;
        pixel_data[75][75] = 0;
        pixel_data[75][76] = 0;
        pixel_data[75][77] = 0;
        pixel_data[75][78] = 0;
        pixel_data[75][79] = 0;
        pixel_data[75][80] = 0;
        pixel_data[75][81] = 0;
        pixel_data[75][82] = 0;
        pixel_data[75][83] = 0;
        pixel_data[75][84] = 0;
        pixel_data[75][85] = 0;
        pixel_data[75][86] = 0;
        pixel_data[75][87] = 0;
        pixel_data[75][88] = 0;
        pixel_data[75][89] = 0;
        pixel_data[75][90] = 0;
        pixel_data[75][91] = 0;
        pixel_data[75][92] = 0;
        pixel_data[75][93] = 0;
        pixel_data[75][94] = 0;
        pixel_data[75][95] = 0;
        pixel_data[75][96] = 0;
        pixel_data[75][97] = 0;
        pixel_data[75][98] = 0;
        pixel_data[75][99] = 0;
        pixel_data[75][100] = 0;
        pixel_data[75][101] = 0;
        pixel_data[75][102] = 0;
        pixel_data[75][103] = 0;
        pixel_data[75][104] = 0;
        pixel_data[75][105] = 0;
        pixel_data[75][106] = 0;
        pixel_data[75][107] = 0;
        pixel_data[75][108] = 0;
        pixel_data[75][109] = 0;
        pixel_data[75][110] = 0;
        pixel_data[75][111] = 0;
        pixel_data[75][112] = 0;
        pixel_data[75][113] = 0;
        pixel_data[75][114] = 0;
        pixel_data[75][115] = 0;
        pixel_data[75][116] = 0;
        pixel_data[75][117] = 0;
        pixel_data[75][118] = 0;
        pixel_data[75][119] = 0;
        pixel_data[75][120] = 0;
        pixel_data[75][121] = 0;
        pixel_data[75][122] = 0;
        pixel_data[75][123] = 0;
        pixel_data[75][124] = 0;
        pixel_data[75][125] = 0;
        pixel_data[75][126] = 0;
        pixel_data[75][127] = 0;
        pixel_data[75][128] = 0;
        pixel_data[75][129] = 0;
        pixel_data[75][130] = 0;
        pixel_data[75][131] = 0;
        pixel_data[75][132] = 0;
        pixel_data[75][133] = 0;
        pixel_data[75][134] = 0;
        pixel_data[75][135] = 0;
        pixel_data[75][136] = 0;
        pixel_data[75][137] = 0;
        pixel_data[75][138] = 0;
        pixel_data[75][139] = 0;
        pixel_data[75][140] = 0;
        pixel_data[75][141] = 0;
        pixel_data[75][142] = 0;
        pixel_data[75][143] = 0;
        pixel_data[75][144] = 0;
        pixel_data[75][145] = 0;
        pixel_data[75][146] = 0;
        pixel_data[75][147] = 0;
        pixel_data[75][148] = 0;
        pixel_data[75][149] = 0;
        pixel_data[75][150] = 0;
        pixel_data[75][151] = 0;
        pixel_data[75][152] = 0;
        pixel_data[75][153] = 0;
        pixel_data[75][154] = 0;
        pixel_data[75][155] = 0;
        pixel_data[75][156] = 0;
        pixel_data[75][157] = 0;
        pixel_data[75][158] = 0;
        pixel_data[75][159] = 0;
        pixel_data[75][160] = 0;
        pixel_data[75][161] = 0;
        pixel_data[75][162] = 0;
        pixel_data[75][163] = 0;
        pixel_data[75][164] = 0;
        pixel_data[75][165] = 0;
        pixel_data[75][166] = 0;
        pixel_data[75][167] = 0;
        pixel_data[75][168] = 0;
        pixel_data[75][169] = 0;
        pixel_data[75][170] = 0;
        pixel_data[75][171] = 0;
        pixel_data[75][172] = 0;
        pixel_data[75][173] = 0;
        pixel_data[75][174] = 0;
        pixel_data[75][175] = 0;
        pixel_data[75][176] = 0;
        pixel_data[75][177] = 0;
        pixel_data[75][178] = 0;
        pixel_data[75][179] = 0;
        pixel_data[75][180] = 0;
        pixel_data[75][181] = 0;
        pixel_data[75][182] = 0;
        pixel_data[75][183] = 0;
        pixel_data[75][184] = 0;
        pixel_data[75][185] = 0;
        pixel_data[75][186] = 0;
        pixel_data[75][187] = 0;
        pixel_data[75][188] = 0;
        pixel_data[75][189] = 0;
        pixel_data[75][190] = 0;
        pixel_data[75][191] = 0;
        pixel_data[75][192] = 0;
        pixel_data[75][193] = 0;
        pixel_data[75][194] = 0;
        pixel_data[75][195] = 0;
        pixel_data[75][196] = 0;
        pixel_data[75][197] = 0;
        pixel_data[75][198] = 0;
        pixel_data[75][199] = 0; // y=75
        pixel_data[76][0] = 0;
        pixel_data[76][1] = 0;
        pixel_data[76][2] = 0;
        pixel_data[76][3] = 0;
        pixel_data[76][4] = 0;
        pixel_data[76][5] = 0;
        pixel_data[76][6] = 0;
        pixel_data[76][7] = 0;
        pixel_data[76][8] = 0;
        pixel_data[76][9] = 0;
        pixel_data[76][10] = 0;
        pixel_data[76][11] = 0;
        pixel_data[76][12] = 0;
        pixel_data[76][13] = 0;
        pixel_data[76][14] = 0;
        pixel_data[76][15] = 0;
        pixel_data[76][16] = 0;
        pixel_data[76][17] = 0;
        pixel_data[76][18] = 0;
        pixel_data[76][19] = 0;
        pixel_data[76][20] = 0;
        pixel_data[76][21] = 0;
        pixel_data[76][22] = 0;
        pixel_data[76][23] = 0;
        pixel_data[76][24] = 0;
        pixel_data[76][25] = 0;
        pixel_data[76][26] = 0;
        pixel_data[76][27] = 0;
        pixel_data[76][28] = 0;
        pixel_data[76][29] = 0;
        pixel_data[76][30] = 0;
        pixel_data[76][31] = 0;
        pixel_data[76][32] = 0;
        pixel_data[76][33] = 0;
        pixel_data[76][34] = 0;
        pixel_data[76][35] = 0;
        pixel_data[76][36] = 0;
        pixel_data[76][37] = 0;
        pixel_data[76][38] = 0;
        pixel_data[76][39] = 0;
        pixel_data[76][40] = 0;
        pixel_data[76][41] = 0;
        pixel_data[76][42] = 0;
        pixel_data[76][43] = 0;
        pixel_data[76][44] = 0;
        pixel_data[76][45] = 0;
        pixel_data[76][46] = 0;
        pixel_data[76][47] = 0;
        pixel_data[76][48] = 0;
        pixel_data[76][49] = 0;
        pixel_data[76][50] = 0;
        pixel_data[76][51] = 0;
        pixel_data[76][52] = 0;
        pixel_data[76][53] = 0;
        pixel_data[76][54] = 0;
        pixel_data[76][55] = 0;
        pixel_data[76][56] = 0;
        pixel_data[76][57] = 0;
        pixel_data[76][58] = 0;
        pixel_data[76][59] = 0;
        pixel_data[76][60] = 0;
        pixel_data[76][61] = 0;
        pixel_data[76][62] = 0;
        pixel_data[76][63] = 0;
        pixel_data[76][64] = 0;
        pixel_data[76][65] = 0;
        pixel_data[76][66] = 0;
        pixel_data[76][67] = 0;
        pixel_data[76][68] = 0;
        pixel_data[76][69] = 0;
        pixel_data[76][70] = 0;
        pixel_data[76][71] = 0;
        pixel_data[76][72] = 0;
        pixel_data[76][73] = 0;
        pixel_data[76][74] = 0;
        pixel_data[76][75] = 0;
        pixel_data[76][76] = 0;
        pixel_data[76][77] = 0;
        pixel_data[76][78] = 0;
        pixel_data[76][79] = 0;
        pixel_data[76][80] = 0;
        pixel_data[76][81] = 0;
        pixel_data[76][82] = 0;
        pixel_data[76][83] = 0;
        pixel_data[76][84] = 0;
        pixel_data[76][85] = 0;
        pixel_data[76][86] = 0;
        pixel_data[76][87] = 0;
        pixel_data[76][88] = 0;
        pixel_data[76][89] = 0;
        pixel_data[76][90] = 0;
        pixel_data[76][91] = 0;
        pixel_data[76][92] = 0;
        pixel_data[76][93] = 0;
        pixel_data[76][94] = 0;
        pixel_data[76][95] = 0;
        pixel_data[76][96] = 0;
        pixel_data[76][97] = 0;
        pixel_data[76][98] = 0;
        pixel_data[76][99] = 0;
        pixel_data[76][100] = 0;
        pixel_data[76][101] = 0;
        pixel_data[76][102] = 0;
        pixel_data[76][103] = 0;
        pixel_data[76][104] = 0;
        pixel_data[76][105] = 0;
        pixel_data[76][106] = 0;
        pixel_data[76][107] = 0;
        pixel_data[76][108] = 0;
        pixel_data[76][109] = 0;
        pixel_data[76][110] = 0;
        pixel_data[76][111] = 0;
        pixel_data[76][112] = 0;
        pixel_data[76][113] = 0;
        pixel_data[76][114] = 0;
        pixel_data[76][115] = 0;
        pixel_data[76][116] = 0;
        pixel_data[76][117] = 0;
        pixel_data[76][118] = 0;
        pixel_data[76][119] = 0;
        pixel_data[76][120] = 0;
        pixel_data[76][121] = 0;
        pixel_data[76][122] = 0;
        pixel_data[76][123] = 0;
        pixel_data[76][124] = 0;
        pixel_data[76][125] = 0;
        pixel_data[76][126] = 0;
        pixel_data[76][127] = 0;
        pixel_data[76][128] = 0;
        pixel_data[76][129] = 0;
        pixel_data[76][130] = 0;
        pixel_data[76][131] = 0;
        pixel_data[76][132] = 0;
        pixel_data[76][133] = 0;
        pixel_data[76][134] = 0;
        pixel_data[76][135] = 0;
        pixel_data[76][136] = 0;
        pixel_data[76][137] = 0;
        pixel_data[76][138] = 0;
        pixel_data[76][139] = 0;
        pixel_data[76][140] = 0;
        pixel_data[76][141] = 0;
        pixel_data[76][142] = 0;
        pixel_data[76][143] = 0;
        pixel_data[76][144] = 0;
        pixel_data[76][145] = 0;
        pixel_data[76][146] = 0;
        pixel_data[76][147] = 0;
        pixel_data[76][148] = 0;
        pixel_data[76][149] = 0;
        pixel_data[76][150] = 0;
        pixel_data[76][151] = 0;
        pixel_data[76][152] = 0;
        pixel_data[76][153] = 0;
        pixel_data[76][154] = 0;
        pixel_data[76][155] = 0;
        pixel_data[76][156] = 0;
        pixel_data[76][157] = 0;
        pixel_data[76][158] = 0;
        pixel_data[76][159] = 0;
        pixel_data[76][160] = 0;
        pixel_data[76][161] = 0;
        pixel_data[76][162] = 0;
        pixel_data[76][163] = 0;
        pixel_data[76][164] = 0;
        pixel_data[76][165] = 0;
        pixel_data[76][166] = 0;
        pixel_data[76][167] = 0;
        pixel_data[76][168] = 0;
        pixel_data[76][169] = 0;
        pixel_data[76][170] = 0;
        pixel_data[76][171] = 0;
        pixel_data[76][172] = 0;
        pixel_data[76][173] = 0;
        pixel_data[76][174] = 0;
        pixel_data[76][175] = 0;
        pixel_data[76][176] = 0;
        pixel_data[76][177] = 0;
        pixel_data[76][178] = 0;
        pixel_data[76][179] = 0;
        pixel_data[76][180] = 0;
        pixel_data[76][181] = 0;
        pixel_data[76][182] = 0;
        pixel_data[76][183] = 0;
        pixel_data[76][184] = 0;
        pixel_data[76][185] = 0;
        pixel_data[76][186] = 0;
        pixel_data[76][187] = 0;
        pixel_data[76][188] = 0;
        pixel_data[76][189] = 0;
        pixel_data[76][190] = 0;
        pixel_data[76][191] = 0;
        pixel_data[76][192] = 0;
        pixel_data[76][193] = 0;
        pixel_data[76][194] = 0;
        pixel_data[76][195] = 0;
        pixel_data[76][196] = 0;
        pixel_data[76][197] = 0;
        pixel_data[76][198] = 0;
        pixel_data[76][199] = 0; // y=76
        pixel_data[77][0] = 0;
        pixel_data[77][1] = 0;
        pixel_data[77][2] = 0;
        pixel_data[77][3] = 0;
        pixel_data[77][4] = 0;
        pixel_data[77][5] = 0;
        pixel_data[77][6] = 0;
        pixel_data[77][7] = 0;
        pixel_data[77][8] = 0;
        pixel_data[77][9] = 0;
        pixel_data[77][10] = 0;
        pixel_data[77][11] = 0;
        pixel_data[77][12] = 0;
        pixel_data[77][13] = 0;
        pixel_data[77][14] = 0;
        pixel_data[77][15] = 0;
        pixel_data[77][16] = 0;
        pixel_data[77][17] = 0;
        pixel_data[77][18] = 0;
        pixel_data[77][19] = 0;
        pixel_data[77][20] = 0;
        pixel_data[77][21] = 0;
        pixel_data[77][22] = 0;
        pixel_data[77][23] = 0;
        pixel_data[77][24] = 0;
        pixel_data[77][25] = 0;
        pixel_data[77][26] = 0;
        pixel_data[77][27] = 0;
        pixel_data[77][28] = 0;
        pixel_data[77][29] = 0;
        pixel_data[77][30] = 0;
        pixel_data[77][31] = 0;
        pixel_data[77][32] = 0;
        pixel_data[77][33] = 0;
        pixel_data[77][34] = 0;
        pixel_data[77][35] = 0;
        pixel_data[77][36] = 0;
        pixel_data[77][37] = 0;
        pixel_data[77][38] = 0;
        pixel_data[77][39] = 0;
        pixel_data[77][40] = 0;
        pixel_data[77][41] = 0;
        pixel_data[77][42] = 0;
        pixel_data[77][43] = 0;
        pixel_data[77][44] = 0;
        pixel_data[77][45] = 0;
        pixel_data[77][46] = 0;
        pixel_data[77][47] = 0;
        pixel_data[77][48] = 0;
        pixel_data[77][49] = 0;
        pixel_data[77][50] = 0;
        pixel_data[77][51] = 0;
        pixel_data[77][52] = 0;
        pixel_data[77][53] = 0;
        pixel_data[77][54] = 0;
        pixel_data[77][55] = 0;
        pixel_data[77][56] = 0;
        pixel_data[77][57] = 0;
        pixel_data[77][58] = 0;
        pixel_data[77][59] = 0;
        pixel_data[77][60] = 0;
        pixel_data[77][61] = 0;
        pixel_data[77][62] = 0;
        pixel_data[77][63] = 0;
        pixel_data[77][64] = 0;
        pixel_data[77][65] = 0;
        pixel_data[77][66] = 0;
        pixel_data[77][67] = 0;
        pixel_data[77][68] = 0;
        pixel_data[77][69] = 0;
        pixel_data[77][70] = 0;
        pixel_data[77][71] = 0;
        pixel_data[77][72] = 0;
        pixel_data[77][73] = 0;
        pixel_data[77][74] = 0;
        pixel_data[77][75] = 0;
        pixel_data[77][76] = 0;
        pixel_data[77][77] = 0;
        pixel_data[77][78] = 0;
        pixel_data[77][79] = 0;
        pixel_data[77][80] = 0;
        pixel_data[77][81] = 0;
        pixel_data[77][82] = 0;
        pixel_data[77][83] = 0;
        pixel_data[77][84] = 0;
        pixel_data[77][85] = 0;
        pixel_data[77][86] = 0;
        pixel_data[77][87] = 0;
        pixel_data[77][88] = 0;
        pixel_data[77][89] = 0;
        pixel_data[77][90] = 0;
        pixel_data[77][91] = 0;
        pixel_data[77][92] = 0;
        pixel_data[77][93] = 0;
        pixel_data[77][94] = 0;
        pixel_data[77][95] = 0;
        pixel_data[77][96] = 0;
        pixel_data[77][97] = 0;
        pixel_data[77][98] = 0;
        pixel_data[77][99] = 0;
        pixel_data[77][100] = 0;
        pixel_data[77][101] = 0;
        pixel_data[77][102] = 0;
        pixel_data[77][103] = 0;
        pixel_data[77][104] = 0;
        pixel_data[77][105] = 0;
        pixel_data[77][106] = 0;
        pixel_data[77][107] = 0;
        pixel_data[77][108] = 0;
        pixel_data[77][109] = 0;
        pixel_data[77][110] = 0;
        pixel_data[77][111] = 0;
        pixel_data[77][112] = 0;
        pixel_data[77][113] = 0;
        pixel_data[77][114] = 0;
        pixel_data[77][115] = 0;
        pixel_data[77][116] = 0;
        pixel_data[77][117] = 0;
        pixel_data[77][118] = 0;
        pixel_data[77][119] = 0;
        pixel_data[77][120] = 0;
        pixel_data[77][121] = 0;
        pixel_data[77][122] = 0;
        pixel_data[77][123] = 0;
        pixel_data[77][124] = 0;
        pixel_data[77][125] = 0;
        pixel_data[77][126] = 0;
        pixel_data[77][127] = 0;
        pixel_data[77][128] = 0;
        pixel_data[77][129] = 0;
        pixel_data[77][130] = 0;
        pixel_data[77][131] = 0;
        pixel_data[77][132] = 0;
        pixel_data[77][133] = 0;
        pixel_data[77][134] = 0;
        pixel_data[77][135] = 0;
        pixel_data[77][136] = 0;
        pixel_data[77][137] = 0;
        pixel_data[77][138] = 0;
        pixel_data[77][139] = 0;
        pixel_data[77][140] = 0;
        pixel_data[77][141] = 0;
        pixel_data[77][142] = 0;
        pixel_data[77][143] = 0;
        pixel_data[77][144] = 0;
        pixel_data[77][145] = 0;
        pixel_data[77][146] = 0;
        pixel_data[77][147] = 0;
        pixel_data[77][148] = 0;
        pixel_data[77][149] = 0;
        pixel_data[77][150] = 0;
        pixel_data[77][151] = 0;
        pixel_data[77][152] = 0;
        pixel_data[77][153] = 0;
        pixel_data[77][154] = 0;
        pixel_data[77][155] = 0;
        pixel_data[77][156] = 0;
        pixel_data[77][157] = 0;
        pixel_data[77][158] = 0;
        pixel_data[77][159] = 0;
        pixel_data[77][160] = 0;
        pixel_data[77][161] = 0;
        pixel_data[77][162] = 0;
        pixel_data[77][163] = 0;
        pixel_data[77][164] = 0;
        pixel_data[77][165] = 0;
        pixel_data[77][166] = 0;
        pixel_data[77][167] = 0;
        pixel_data[77][168] = 0;
        pixel_data[77][169] = 0;
        pixel_data[77][170] = 0;
        pixel_data[77][171] = 0;
        pixel_data[77][172] = 0;
        pixel_data[77][173] = 0;
        pixel_data[77][174] = 0;
        pixel_data[77][175] = 0;
        pixel_data[77][176] = 0;
        pixel_data[77][177] = 0;
        pixel_data[77][178] = 0;
        pixel_data[77][179] = 0;
        pixel_data[77][180] = 0;
        pixel_data[77][181] = 0;
        pixel_data[77][182] = 0;
        pixel_data[77][183] = 0;
        pixel_data[77][184] = 0;
        pixel_data[77][185] = 0;
        pixel_data[77][186] = 0;
        pixel_data[77][187] = 0;
        pixel_data[77][188] = 0;
        pixel_data[77][189] = 0;
        pixel_data[77][190] = 0;
        pixel_data[77][191] = 0;
        pixel_data[77][192] = 0;
        pixel_data[77][193] = 0;
        pixel_data[77][194] = 0;
        pixel_data[77][195] = 0;
        pixel_data[77][196] = 0;
        pixel_data[77][197] = 0;
        pixel_data[77][198] = 0;
        pixel_data[77][199] = 0; // y=77
        pixel_data[78][0] = 0;
        pixel_data[78][1] = 0;
        pixel_data[78][2] = 0;
        pixel_data[78][3] = 0;
        pixel_data[78][4] = 0;
        pixel_data[78][5] = 0;
        pixel_data[78][6] = 0;
        pixel_data[78][7] = 0;
        pixel_data[78][8] = 0;
        pixel_data[78][9] = 0;
        pixel_data[78][10] = 0;
        pixel_data[78][11] = 0;
        pixel_data[78][12] = 0;
        pixel_data[78][13] = 0;
        pixel_data[78][14] = 0;
        pixel_data[78][15] = 0;
        pixel_data[78][16] = 0;
        pixel_data[78][17] = 0;
        pixel_data[78][18] = 0;
        pixel_data[78][19] = 0;
        pixel_data[78][20] = 0;
        pixel_data[78][21] = 0;
        pixel_data[78][22] = 0;
        pixel_data[78][23] = 0;
        pixel_data[78][24] = 0;
        pixel_data[78][25] = 0;
        pixel_data[78][26] = 0;
        pixel_data[78][27] = 0;
        pixel_data[78][28] = 0;
        pixel_data[78][29] = 0;
        pixel_data[78][30] = 0;
        pixel_data[78][31] = 0;
        pixel_data[78][32] = 0;
        pixel_data[78][33] = 0;
        pixel_data[78][34] = 0;
        pixel_data[78][35] = 0;
        pixel_data[78][36] = 0;
        pixel_data[78][37] = 0;
        pixel_data[78][38] = 0;
        pixel_data[78][39] = 0;
        pixel_data[78][40] = 0;
        pixel_data[78][41] = 0;
        pixel_data[78][42] = 0;
        pixel_data[78][43] = 0;
        pixel_data[78][44] = 0;
        pixel_data[78][45] = 0;
        pixel_data[78][46] = 0;
        pixel_data[78][47] = 0;
        pixel_data[78][48] = 0;
        pixel_data[78][49] = 0;
        pixel_data[78][50] = 0;
        pixel_data[78][51] = 0;
        pixel_data[78][52] = 0;
        pixel_data[78][53] = 0;
        pixel_data[78][54] = 0;
        pixel_data[78][55] = 0;
        pixel_data[78][56] = 0;
        pixel_data[78][57] = 0;
        pixel_data[78][58] = 0;
        pixel_data[78][59] = 0;
        pixel_data[78][60] = 0;
        pixel_data[78][61] = 0;
        pixel_data[78][62] = 0;
        pixel_data[78][63] = 0;
        pixel_data[78][64] = 0;
        pixel_data[78][65] = 0;
        pixel_data[78][66] = 0;
        pixel_data[78][67] = 0;
        pixel_data[78][68] = 0;
        pixel_data[78][69] = 0;
        pixel_data[78][70] = 0;
        pixel_data[78][71] = 0;
        pixel_data[78][72] = 0;
        pixel_data[78][73] = 0;
        pixel_data[78][74] = 0;
        pixel_data[78][75] = 0;
        pixel_data[78][76] = 0;
        pixel_data[78][77] = 0;
        pixel_data[78][78] = 0;
        pixel_data[78][79] = 0;
        pixel_data[78][80] = 0;
        pixel_data[78][81] = 0;
        pixel_data[78][82] = 0;
        pixel_data[78][83] = 0;
        pixel_data[78][84] = 0;
        pixel_data[78][85] = 0;
        pixel_data[78][86] = 0;
        pixel_data[78][87] = 0;
        pixel_data[78][88] = 0;
        pixel_data[78][89] = 0;
        pixel_data[78][90] = 0;
        pixel_data[78][91] = 0;
        pixel_data[78][92] = 0;
        pixel_data[78][93] = 0;
        pixel_data[78][94] = 0;
        pixel_data[78][95] = 0;
        pixel_data[78][96] = 0;
        pixel_data[78][97] = 0;
        pixel_data[78][98] = 0;
        pixel_data[78][99] = 0;
        pixel_data[78][100] = 0;
        pixel_data[78][101] = 0;
        pixel_data[78][102] = 0;
        pixel_data[78][103] = 0;
        pixel_data[78][104] = 0;
        pixel_data[78][105] = 0;
        pixel_data[78][106] = 0;
        pixel_data[78][107] = 0;
        pixel_data[78][108] = 0;
        pixel_data[78][109] = 0;
        pixel_data[78][110] = 0;
        pixel_data[78][111] = 0;
        pixel_data[78][112] = 0;
        pixel_data[78][113] = 0;
        pixel_data[78][114] = 0;
        pixel_data[78][115] = 0;
        pixel_data[78][116] = 0;
        pixel_data[78][117] = 0;
        pixel_data[78][118] = 0;
        pixel_data[78][119] = 0;
        pixel_data[78][120] = 0;
        pixel_data[78][121] = 0;
        pixel_data[78][122] = 0;
        pixel_data[78][123] = 0;
        pixel_data[78][124] = 0;
        pixel_data[78][125] = 0;
        pixel_data[78][126] = 0;
        pixel_data[78][127] = 0;
        pixel_data[78][128] = 0;
        pixel_data[78][129] = 0;
        pixel_data[78][130] = 0;
        pixel_data[78][131] = 0;
        pixel_data[78][132] = 0;
        pixel_data[78][133] = 0;
        pixel_data[78][134] = 0;
        pixel_data[78][135] = 0;
        pixel_data[78][136] = 0;
        pixel_data[78][137] = 0;
        pixel_data[78][138] = 0;
        pixel_data[78][139] = 0;
        pixel_data[78][140] = 0;
        pixel_data[78][141] = 0;
        pixel_data[78][142] = 0;
        pixel_data[78][143] = 0;
        pixel_data[78][144] = 0;
        pixel_data[78][145] = 0;
        pixel_data[78][146] = 0;
        pixel_data[78][147] = 0;
        pixel_data[78][148] = 0;
        pixel_data[78][149] = 0;
        pixel_data[78][150] = 0;
        pixel_data[78][151] = 0;
        pixel_data[78][152] = 0;
        pixel_data[78][153] = 0;
        pixel_data[78][154] = 0;
        pixel_data[78][155] = 0;
        pixel_data[78][156] = 0;
        pixel_data[78][157] = 0;
        pixel_data[78][158] = 0;
        pixel_data[78][159] = 0;
        pixel_data[78][160] = 0;
        pixel_data[78][161] = 0;
        pixel_data[78][162] = 0;
        pixel_data[78][163] = 0;
        pixel_data[78][164] = 0;
        pixel_data[78][165] = 0;
        pixel_data[78][166] = 0;
        pixel_data[78][167] = 0;
        pixel_data[78][168] = 0;
        pixel_data[78][169] = 0;
        pixel_data[78][170] = 0;
        pixel_data[78][171] = 0;
        pixel_data[78][172] = 0;
        pixel_data[78][173] = 0;
        pixel_data[78][174] = 0;
        pixel_data[78][175] = 0;
        pixel_data[78][176] = 0;
        pixel_data[78][177] = 0;
        pixel_data[78][178] = 0;
        pixel_data[78][179] = 0;
        pixel_data[78][180] = 0;
        pixel_data[78][181] = 0;
        pixel_data[78][182] = 0;
        pixel_data[78][183] = 0;
        pixel_data[78][184] = 0;
        pixel_data[78][185] = 0;
        pixel_data[78][186] = 0;
        pixel_data[78][187] = 0;
        pixel_data[78][188] = 0;
        pixel_data[78][189] = 0;
        pixel_data[78][190] = 0;
        pixel_data[78][191] = 0;
        pixel_data[78][192] = 0;
        pixel_data[78][193] = 0;
        pixel_data[78][194] = 0;
        pixel_data[78][195] = 0;
        pixel_data[78][196] = 0;
        pixel_data[78][197] = 0;
        pixel_data[78][198] = 0;
        pixel_data[78][199] = 0; // y=78
        pixel_data[79][0] = 0;
        pixel_data[79][1] = 0;
        pixel_data[79][2] = 0;
        pixel_data[79][3] = 0;
        pixel_data[79][4] = 0;
        pixel_data[79][5] = 0;
        pixel_data[79][6] = 0;
        pixel_data[79][7] = 0;
        pixel_data[79][8] = 0;
        pixel_data[79][9] = 0;
        pixel_data[79][10] = 0;
        pixel_data[79][11] = 0;
        pixel_data[79][12] = 0;
        pixel_data[79][13] = 0;
        pixel_data[79][14] = 0;
        pixel_data[79][15] = 0;
        pixel_data[79][16] = 0;
        pixel_data[79][17] = 0;
        pixel_data[79][18] = 0;
        pixel_data[79][19] = 0;
        pixel_data[79][20] = 0;
        pixel_data[79][21] = 0;
        pixel_data[79][22] = 0;
        pixel_data[79][23] = 0;
        pixel_data[79][24] = 0;
        pixel_data[79][25] = 0;
        pixel_data[79][26] = 0;
        pixel_data[79][27] = 0;
        pixel_data[79][28] = 0;
        pixel_data[79][29] = 0;
        pixel_data[79][30] = 0;
        pixel_data[79][31] = 0;
        pixel_data[79][32] = 0;
        pixel_data[79][33] = 0;
        pixel_data[79][34] = 0;
        pixel_data[79][35] = 0;
        pixel_data[79][36] = 0;
        pixel_data[79][37] = 0;
        pixel_data[79][38] = 0;
        pixel_data[79][39] = 0;
        pixel_data[79][40] = 0;
        pixel_data[79][41] = 0;
        pixel_data[79][42] = 0;
        pixel_data[79][43] = 0;
        pixel_data[79][44] = 0;
        pixel_data[79][45] = 0;
        pixel_data[79][46] = 0;
        pixel_data[79][47] = 0;
        pixel_data[79][48] = 0;
        pixel_data[79][49] = 0;
        pixel_data[79][50] = 0;
        pixel_data[79][51] = 0;
        pixel_data[79][52] = 0;
        pixel_data[79][53] = 0;
        pixel_data[79][54] = 0;
        pixel_data[79][55] = 0;
        pixel_data[79][56] = 0;
        pixel_data[79][57] = 0;
        pixel_data[79][58] = 0;
        pixel_data[79][59] = 0;
        pixel_data[79][60] = 0;
        pixel_data[79][61] = 0;
        pixel_data[79][62] = 0;
        pixel_data[79][63] = 0;
        pixel_data[79][64] = 0;
        pixel_data[79][65] = 0;
        pixel_data[79][66] = 0;
        pixel_data[79][67] = 0;
        pixel_data[79][68] = 0;
        pixel_data[79][69] = 0;
        pixel_data[79][70] = 0;
        pixel_data[79][71] = 0;
        pixel_data[79][72] = 0;
        pixel_data[79][73] = 0;
        pixel_data[79][74] = 0;
        pixel_data[79][75] = 0;
        pixel_data[79][76] = 0;
        pixel_data[79][77] = 0;
        pixel_data[79][78] = 0;
        pixel_data[79][79] = 0;
        pixel_data[79][80] = 0;
        pixel_data[79][81] = 0;
        pixel_data[79][82] = 0;
        pixel_data[79][83] = 0;
        pixel_data[79][84] = 0;
        pixel_data[79][85] = 0;
        pixel_data[79][86] = 0;
        pixel_data[79][87] = 0;
        pixel_data[79][88] = 0;
        pixel_data[79][89] = 0;
        pixel_data[79][90] = 0;
        pixel_data[79][91] = 0;
        pixel_data[79][92] = 0;
        pixel_data[79][93] = 0;
        pixel_data[79][94] = 0;
        pixel_data[79][95] = 0;
        pixel_data[79][96] = 0;
        pixel_data[79][97] = 0;
        pixel_data[79][98] = 0;
        pixel_data[79][99] = 0;
        pixel_data[79][100] = 0;
        pixel_data[79][101] = 0;
        pixel_data[79][102] = 0;
        pixel_data[79][103] = 0;
        pixel_data[79][104] = 0;
        pixel_data[79][105] = 0;
        pixel_data[79][106] = 0;
        pixel_data[79][107] = 0;
        pixel_data[79][108] = 0;
        pixel_data[79][109] = 0;
        pixel_data[79][110] = 0;
        pixel_data[79][111] = 0;
        pixel_data[79][112] = 0;
        pixel_data[79][113] = 0;
        pixel_data[79][114] = 0;
        pixel_data[79][115] = 0;
        pixel_data[79][116] = 0;
        pixel_data[79][117] = 0;
        pixel_data[79][118] = 0;
        pixel_data[79][119] = 0;
        pixel_data[79][120] = 0;
        pixel_data[79][121] = 0;
        pixel_data[79][122] = 0;
        pixel_data[79][123] = 0;
        pixel_data[79][124] = 0;
        pixel_data[79][125] = 0;
        pixel_data[79][126] = 0;
        pixel_data[79][127] = 0;
        pixel_data[79][128] = 0;
        pixel_data[79][129] = 0;
        pixel_data[79][130] = 0;
        pixel_data[79][131] = 0;
        pixel_data[79][132] = 0;
        pixel_data[79][133] = 0;
        pixel_data[79][134] = 0;
        pixel_data[79][135] = 0;
        pixel_data[79][136] = 0;
        pixel_data[79][137] = 0;
        pixel_data[79][138] = 0;
        pixel_data[79][139] = 0;
        pixel_data[79][140] = 0;
        pixel_data[79][141] = 0;
        pixel_data[79][142] = 0;
        pixel_data[79][143] = 0;
        pixel_data[79][144] = 0;
        pixel_data[79][145] = 0;
        pixel_data[79][146] = 0;
        pixel_data[79][147] = 0;
        pixel_data[79][148] = 0;
        pixel_data[79][149] = 0;
        pixel_data[79][150] = 0;
        pixel_data[79][151] = 0;
        pixel_data[79][152] = 0;
        pixel_data[79][153] = 0;
        pixel_data[79][154] = 0;
        pixel_data[79][155] = 0;
        pixel_data[79][156] = 0;
        pixel_data[79][157] = 0;
        pixel_data[79][158] = 0;
        pixel_data[79][159] = 0;
        pixel_data[79][160] = 0;
        pixel_data[79][161] = 0;
        pixel_data[79][162] = 0;
        pixel_data[79][163] = 0;
        pixel_data[79][164] = 0;
        pixel_data[79][165] = 0;
        pixel_data[79][166] = 0;
        pixel_data[79][167] = 0;
        pixel_data[79][168] = 0;
        pixel_data[79][169] = 0;
        pixel_data[79][170] = 0;
        pixel_data[79][171] = 0;
        pixel_data[79][172] = 0;
        pixel_data[79][173] = 0;
        pixel_data[79][174] = 0;
        pixel_data[79][175] = 0;
        pixel_data[79][176] = 0;
        pixel_data[79][177] = 0;
        pixel_data[79][178] = 0;
        pixel_data[79][179] = 0;
        pixel_data[79][180] = 0;
        pixel_data[79][181] = 0;
        pixel_data[79][182] = 0;
        pixel_data[79][183] = 0;
        pixel_data[79][184] = 0;
        pixel_data[79][185] = 0;
        pixel_data[79][186] = 0;
        pixel_data[79][187] = 0;
        pixel_data[79][188] = 0;
        pixel_data[79][189] = 0;
        pixel_data[79][190] = 0;
        pixel_data[79][191] = 0;
        pixel_data[79][192] = 0;
        pixel_data[79][193] = 0;
        pixel_data[79][194] = 0;
        pixel_data[79][195] = 0;
        pixel_data[79][196] = 0;
        pixel_data[79][197] = 0;
        pixel_data[79][198] = 0;
        pixel_data[79][199] = 0; // y=79
        pixel_data[80][0] = 0;
        pixel_data[80][1] = 0;
        pixel_data[80][2] = 0;
        pixel_data[80][3] = 0;
        pixel_data[80][4] = 0;
        pixel_data[80][5] = 0;
        pixel_data[80][6] = 0;
        pixel_data[80][7] = 0;
        pixel_data[80][8] = 0;
        pixel_data[80][9] = 0;
        pixel_data[80][10] = 0;
        pixel_data[80][11] = 0;
        pixel_data[80][12] = 0;
        pixel_data[80][13] = 0;
        pixel_data[80][14] = 0;
        pixel_data[80][15] = 0;
        pixel_data[80][16] = 0;
        pixel_data[80][17] = 0;
        pixel_data[80][18] = 0;
        pixel_data[80][19] = 0;
        pixel_data[80][20] = 0;
        pixel_data[80][21] = 0;
        pixel_data[80][22] = 0;
        pixel_data[80][23] = 0;
        pixel_data[80][24] = 0;
        pixel_data[80][25] = 0;
        pixel_data[80][26] = 0;
        pixel_data[80][27] = 0;
        pixel_data[80][28] = 0;
        pixel_data[80][29] = 0;
        pixel_data[80][30] = 0;
        pixel_data[80][31] = 0;
        pixel_data[80][32] = 0;
        pixel_data[80][33] = 0;
        pixel_data[80][34] = 0;
        pixel_data[80][35] = 0;
        pixel_data[80][36] = 0;
        pixel_data[80][37] = 0;
        pixel_data[80][38] = 0;
        pixel_data[80][39] = 0;
        pixel_data[80][40] = 0;
        pixel_data[80][41] = 0;
        pixel_data[80][42] = 0;
        pixel_data[80][43] = 0;
        pixel_data[80][44] = 0;
        pixel_data[80][45] = 0;
        pixel_data[80][46] = 0;
        pixel_data[80][47] = 0;
        pixel_data[80][48] = 0;
        pixel_data[80][49] = 0;
        pixel_data[80][50] = 0;
        pixel_data[80][51] = 0;
        pixel_data[80][52] = 0;
        pixel_data[80][53] = 0;
        pixel_data[80][54] = 0;
        pixel_data[80][55] = 0;
        pixel_data[80][56] = 0;
        pixel_data[80][57] = 0;
        pixel_data[80][58] = 0;
        pixel_data[80][59] = 0;
        pixel_data[80][60] = 0;
        pixel_data[80][61] = 0;
        pixel_data[80][62] = 0;
        pixel_data[80][63] = 0;
        pixel_data[80][64] = 0;
        pixel_data[80][65] = 0;
        pixel_data[80][66] = 0;
        pixel_data[80][67] = 0;
        pixel_data[80][68] = 0;
        pixel_data[80][69] = 0;
        pixel_data[80][70] = 0;
        pixel_data[80][71] = 0;
        pixel_data[80][72] = 0;
        pixel_data[80][73] = 0;
        pixel_data[80][74] = 0;
        pixel_data[80][75] = 0;
        pixel_data[80][76] = 0;
        pixel_data[80][77] = 0;
        pixel_data[80][78] = 0;
        pixel_data[80][79] = 0;
        pixel_data[80][80] = 0;
        pixel_data[80][81] = 0;
        pixel_data[80][82] = 0;
        pixel_data[80][83] = 0;
        pixel_data[80][84] = 0;
        pixel_data[80][85] = 0;
        pixel_data[80][86] = 0;
        pixel_data[80][87] = 0;
        pixel_data[80][88] = 0;
        pixel_data[80][89] = 0;
        pixel_data[80][90] = 0;
        pixel_data[80][91] = 0;
        pixel_data[80][92] = 0;
        pixel_data[80][93] = 0;
        pixel_data[80][94] = 0;
        pixel_data[80][95] = 0;
        pixel_data[80][96] = 0;
        pixel_data[80][97] = 0;
        pixel_data[80][98] = 0;
        pixel_data[80][99] = 0;
        pixel_data[80][100] = 0;
        pixel_data[80][101] = 0;
        pixel_data[80][102] = 0;
        pixel_data[80][103] = 0;
        pixel_data[80][104] = 0;
        pixel_data[80][105] = 0;
        pixel_data[80][106] = 0;
        pixel_data[80][107] = 0;
        pixel_data[80][108] = 0;
        pixel_data[80][109] = 0;
        pixel_data[80][110] = 0;
        pixel_data[80][111] = 0;
        pixel_data[80][112] = 0;
        pixel_data[80][113] = 0;
        pixel_data[80][114] = 0;
        pixel_data[80][115] = 0;
        pixel_data[80][116] = 0;
        pixel_data[80][117] = 0;
        pixel_data[80][118] = 0;
        pixel_data[80][119] = 0;
        pixel_data[80][120] = 0;
        pixel_data[80][121] = 0;
        pixel_data[80][122] = 0;
        pixel_data[80][123] = 0;
        pixel_data[80][124] = 0;
        pixel_data[80][125] = 0;
        pixel_data[80][126] = 0;
        pixel_data[80][127] = 0;
        pixel_data[80][128] = 0;
        pixel_data[80][129] = 0;
        pixel_data[80][130] = 0;
        pixel_data[80][131] = 0;
        pixel_data[80][132] = 0;
        pixel_data[80][133] = 0;
        pixel_data[80][134] = 0;
        pixel_data[80][135] = 0;
        pixel_data[80][136] = 0;
        pixel_data[80][137] = 0;
        pixel_data[80][138] = 0;
        pixel_data[80][139] = 0;
        pixel_data[80][140] = 0;
        pixel_data[80][141] = 0;
        pixel_data[80][142] = 0;
        pixel_data[80][143] = 0;
        pixel_data[80][144] = 0;
        pixel_data[80][145] = 0;
        pixel_data[80][146] = 0;
        pixel_data[80][147] = 0;
        pixel_data[80][148] = 0;
        pixel_data[80][149] = 0;
        pixel_data[80][150] = 0;
        pixel_data[80][151] = 0;
        pixel_data[80][152] = 0;
        pixel_data[80][153] = 0;
        pixel_data[80][154] = 0;
        pixel_data[80][155] = 0;
        pixel_data[80][156] = 0;
        pixel_data[80][157] = 0;
        pixel_data[80][158] = 0;
        pixel_data[80][159] = 0;
        pixel_data[80][160] = 0;
        pixel_data[80][161] = 0;
        pixel_data[80][162] = 0;
        pixel_data[80][163] = 0;
        pixel_data[80][164] = 0;
        pixel_data[80][165] = 0;
        pixel_data[80][166] = 0;
        pixel_data[80][167] = 0;
        pixel_data[80][168] = 0;
        pixel_data[80][169] = 0;
        pixel_data[80][170] = 0;
        pixel_data[80][171] = 0;
        pixel_data[80][172] = 0;
        pixel_data[80][173] = 0;
        pixel_data[80][174] = 0;
        pixel_data[80][175] = 0;
        pixel_data[80][176] = 0;
        pixel_data[80][177] = 0;
        pixel_data[80][178] = 0;
        pixel_data[80][179] = 0;
        pixel_data[80][180] = 0;
        pixel_data[80][181] = 0;
        pixel_data[80][182] = 0;
        pixel_data[80][183] = 0;
        pixel_data[80][184] = 0;
        pixel_data[80][185] = 0;
        pixel_data[80][186] = 0;
        pixel_data[80][187] = 0;
        pixel_data[80][188] = 0;
        pixel_data[80][189] = 0;
        pixel_data[80][190] = 0;
        pixel_data[80][191] = 0;
        pixel_data[80][192] = 0;
        pixel_data[80][193] = 0;
        pixel_data[80][194] = 0;
        pixel_data[80][195] = 0;
        pixel_data[80][196] = 0;
        pixel_data[80][197] = 0;
        pixel_data[80][198] = 0;
        pixel_data[80][199] = 0; // y=80
        pixel_data[81][0] = 0;
        pixel_data[81][1] = 0;
        pixel_data[81][2] = 0;
        pixel_data[81][3] = 0;
        pixel_data[81][4] = 0;
        pixel_data[81][5] = 0;
        pixel_data[81][6] = 0;
        pixel_data[81][7] = 0;
        pixel_data[81][8] = 0;
        pixel_data[81][9] = 0;
        pixel_data[81][10] = 0;
        pixel_data[81][11] = 0;
        pixel_data[81][12] = 0;
        pixel_data[81][13] = 0;
        pixel_data[81][14] = 0;
        pixel_data[81][15] = 0;
        pixel_data[81][16] = 0;
        pixel_data[81][17] = 0;
        pixel_data[81][18] = 0;
        pixel_data[81][19] = 0;
        pixel_data[81][20] = 0;
        pixel_data[81][21] = 0;
        pixel_data[81][22] = 0;
        pixel_data[81][23] = 0;
        pixel_data[81][24] = 0;
        pixel_data[81][25] = 0;
        pixel_data[81][26] = 0;
        pixel_data[81][27] = 0;
        pixel_data[81][28] = 0;
        pixel_data[81][29] = 0;
        pixel_data[81][30] = 0;
        pixel_data[81][31] = 0;
        pixel_data[81][32] = 0;
        pixel_data[81][33] = 0;
        pixel_data[81][34] = 0;
        pixel_data[81][35] = 0;
        pixel_data[81][36] = 0;
        pixel_data[81][37] = 0;
        pixel_data[81][38] = 0;
        pixel_data[81][39] = 0;
        pixel_data[81][40] = 0;
        pixel_data[81][41] = 0;
        pixel_data[81][42] = 0;
        pixel_data[81][43] = 0;
        pixel_data[81][44] = 0;
        pixel_data[81][45] = 0;
        pixel_data[81][46] = 0;
        pixel_data[81][47] = 0;
        pixel_data[81][48] = 0;
        pixel_data[81][49] = 0;
        pixel_data[81][50] = 0;
        pixel_data[81][51] = 0;
        pixel_data[81][52] = 0;
        pixel_data[81][53] = 0;
        pixel_data[81][54] = 0;
        pixel_data[81][55] = 0;
        pixel_data[81][56] = 0;
        pixel_data[81][57] = 0;
        pixel_data[81][58] = 0;
        pixel_data[81][59] = 0;
        pixel_data[81][60] = 0;
        pixel_data[81][61] = 0;
        pixel_data[81][62] = 0;
        pixel_data[81][63] = 0;
        pixel_data[81][64] = 0;
        pixel_data[81][65] = 0;
        pixel_data[81][66] = 0;
        pixel_data[81][67] = 0;
        pixel_data[81][68] = 0;
        pixel_data[81][69] = 0;
        pixel_data[81][70] = 0;
        pixel_data[81][71] = 0;
        pixel_data[81][72] = 0;
        pixel_data[81][73] = 0;
        pixel_data[81][74] = 0;
        pixel_data[81][75] = 0;
        pixel_data[81][76] = 0;
        pixel_data[81][77] = 0;
        pixel_data[81][78] = 0;
        pixel_data[81][79] = 0;
        pixel_data[81][80] = 0;
        pixel_data[81][81] = 0;
        pixel_data[81][82] = 0;
        pixel_data[81][83] = 0;
        pixel_data[81][84] = 0;
        pixel_data[81][85] = 0;
        pixel_data[81][86] = 0;
        pixel_data[81][87] = 0;
        pixel_data[81][88] = 0;
        pixel_data[81][89] = 0;
        pixel_data[81][90] = 0;
        pixel_data[81][91] = 0;
        pixel_data[81][92] = 0;
        pixel_data[81][93] = 0;
        pixel_data[81][94] = 0;
        pixel_data[81][95] = 0;
        pixel_data[81][96] = 0;
        pixel_data[81][97] = 0;
        pixel_data[81][98] = 0;
        pixel_data[81][99] = 0;
        pixel_data[81][100] = 0;
        pixel_data[81][101] = 0;
        pixel_data[81][102] = 0;
        pixel_data[81][103] = 0;
        pixel_data[81][104] = 0;
        pixel_data[81][105] = 0;
        pixel_data[81][106] = 0;
        pixel_data[81][107] = 0;
        pixel_data[81][108] = 0;
        pixel_data[81][109] = 0;
        pixel_data[81][110] = 0;
        pixel_data[81][111] = 0;
        pixel_data[81][112] = 0;
        pixel_data[81][113] = 0;
        pixel_data[81][114] = 0;
        pixel_data[81][115] = 0;
        pixel_data[81][116] = 0;
        pixel_data[81][117] = 0;
        pixel_data[81][118] = 0;
        pixel_data[81][119] = 0;
        pixel_data[81][120] = 0;
        pixel_data[81][121] = 0;
        pixel_data[81][122] = 0;
        pixel_data[81][123] = 0;
        pixel_data[81][124] = 0;
        pixel_data[81][125] = 0;
        pixel_data[81][126] = 0;
        pixel_data[81][127] = 0;
        pixel_data[81][128] = 0;
        pixel_data[81][129] = 0;
        pixel_data[81][130] = 0;
        pixel_data[81][131] = 0;
        pixel_data[81][132] = 0;
        pixel_data[81][133] = 0;
        pixel_data[81][134] = 0;
        pixel_data[81][135] = 0;
        pixel_data[81][136] = 0;
        pixel_data[81][137] = 0;
        pixel_data[81][138] = 0;
        pixel_data[81][139] = 0;
        pixel_data[81][140] = 0;
        pixel_data[81][141] = 0;
        pixel_data[81][142] = 0;
        pixel_data[81][143] = 0;
        pixel_data[81][144] = 0;
        pixel_data[81][145] = 0;
        pixel_data[81][146] = 0;
        pixel_data[81][147] = 0;
        pixel_data[81][148] = 0;
        pixel_data[81][149] = 0;
        pixel_data[81][150] = 0;
        pixel_data[81][151] = 0;
        pixel_data[81][152] = 0;
        pixel_data[81][153] = 0;
        pixel_data[81][154] = 0;
        pixel_data[81][155] = 0;
        pixel_data[81][156] = 0;
        pixel_data[81][157] = 0;
        pixel_data[81][158] = 0;
        pixel_data[81][159] = 0;
        pixel_data[81][160] = 0;
        pixel_data[81][161] = 0;
        pixel_data[81][162] = 0;
        pixel_data[81][163] = 0;
        pixel_data[81][164] = 0;
        pixel_data[81][165] = 0;
        pixel_data[81][166] = 0;
        pixel_data[81][167] = 0;
        pixel_data[81][168] = 0;
        pixel_data[81][169] = 0;
        pixel_data[81][170] = 0;
        pixel_data[81][171] = 0;
        pixel_data[81][172] = 0;
        pixel_data[81][173] = 0;
        pixel_data[81][174] = 0;
        pixel_data[81][175] = 0;
        pixel_data[81][176] = 0;
        pixel_data[81][177] = 0;
        pixel_data[81][178] = 0;
        pixel_data[81][179] = 0;
        pixel_data[81][180] = 0;
        pixel_data[81][181] = 0;
        pixel_data[81][182] = 0;
        pixel_data[81][183] = 0;
        pixel_data[81][184] = 0;
        pixel_data[81][185] = 0;
        pixel_data[81][186] = 0;
        pixel_data[81][187] = 0;
        pixel_data[81][188] = 0;
        pixel_data[81][189] = 0;
        pixel_data[81][190] = 0;
        pixel_data[81][191] = 0;
        pixel_data[81][192] = 0;
        pixel_data[81][193] = 0;
        pixel_data[81][194] = 0;
        pixel_data[81][195] = 0;
        pixel_data[81][196] = 0;
        pixel_data[81][197] = 0;
        pixel_data[81][198] = 0;
        pixel_data[81][199] = 0; // y=81
        pixel_data[82][0] = 0;
        pixel_data[82][1] = 0;
        pixel_data[82][2] = 0;
        pixel_data[82][3] = 0;
        pixel_data[82][4] = 0;
        pixel_data[82][5] = 0;
        pixel_data[82][6] = 0;
        pixel_data[82][7] = 0;
        pixel_data[82][8] = 0;
        pixel_data[82][9] = 0;
        pixel_data[82][10] = 0;
        pixel_data[82][11] = 0;
        pixel_data[82][12] = 0;
        pixel_data[82][13] = 0;
        pixel_data[82][14] = 0;
        pixel_data[82][15] = 0;
        pixel_data[82][16] = 0;
        pixel_data[82][17] = 0;
        pixel_data[82][18] = 0;
        pixel_data[82][19] = 0;
        pixel_data[82][20] = 0;
        pixel_data[82][21] = 0;
        pixel_data[82][22] = 0;
        pixel_data[82][23] = 0;
        pixel_data[82][24] = 0;
        pixel_data[82][25] = 0;
        pixel_data[82][26] = 0;
        pixel_data[82][27] = 0;
        pixel_data[82][28] = 0;
        pixel_data[82][29] = 0;
        pixel_data[82][30] = 0;
        pixel_data[82][31] = 0;
        pixel_data[82][32] = 0;
        pixel_data[82][33] = 0;
        pixel_data[82][34] = 0;
        pixel_data[82][35] = 0;
        pixel_data[82][36] = 0;
        pixel_data[82][37] = 0;
        pixel_data[82][38] = 0;
        pixel_data[82][39] = 0;
        pixel_data[82][40] = 0;
        pixel_data[82][41] = 0;
        pixel_data[82][42] = 0;
        pixel_data[82][43] = 0;
        pixel_data[82][44] = 0;
        pixel_data[82][45] = 0;
        pixel_data[82][46] = 0;
        pixel_data[82][47] = 0;
        pixel_data[82][48] = 0;
        pixel_data[82][49] = 0;
        pixel_data[82][50] = 0;
        pixel_data[82][51] = 0;
        pixel_data[82][52] = 0;
        pixel_data[82][53] = 0;
        pixel_data[82][54] = 0;
        pixel_data[82][55] = 0;
        pixel_data[82][56] = 0;
        pixel_data[82][57] = 0;
        pixel_data[82][58] = 0;
        pixel_data[82][59] = 0;
        pixel_data[82][60] = 0;
        pixel_data[82][61] = 0;
        pixel_data[82][62] = 0;
        pixel_data[82][63] = 0;
        pixel_data[82][64] = 0;
        pixel_data[82][65] = 0;
        pixel_data[82][66] = 0;
        pixel_data[82][67] = 0;
        pixel_data[82][68] = 0;
        pixel_data[82][69] = 0;
        pixel_data[82][70] = 0;
        pixel_data[82][71] = 0;
        pixel_data[82][72] = 0;
        pixel_data[82][73] = 0;
        pixel_data[82][74] = 0;
        pixel_data[82][75] = 0;
        pixel_data[82][76] = 0;
        pixel_data[82][77] = 0;
        pixel_data[82][78] = 0;
        pixel_data[82][79] = 0;
        pixel_data[82][80] = 0;
        pixel_data[82][81] = 0;
        pixel_data[82][82] = 0;
        pixel_data[82][83] = 0;
        pixel_data[82][84] = 0;
        pixel_data[82][85] = 0;
        pixel_data[82][86] = 0;
        pixel_data[82][87] = 0;
        pixel_data[82][88] = 0;
        pixel_data[82][89] = 0;
        pixel_data[82][90] = 0;
        pixel_data[82][91] = 0;
        pixel_data[82][92] = 0;
        pixel_data[82][93] = 0;
        pixel_data[82][94] = 0;
        pixel_data[82][95] = 0;
        pixel_data[82][96] = 0;
        pixel_data[82][97] = 0;
        pixel_data[82][98] = 0;
        pixel_data[82][99] = 0;
        pixel_data[82][100] = 0;
        pixel_data[82][101] = 0;
        pixel_data[82][102] = 0;
        pixel_data[82][103] = 0;
        pixel_data[82][104] = 0;
        pixel_data[82][105] = 0;
        pixel_data[82][106] = 0;
        pixel_data[82][107] = 0;
        pixel_data[82][108] = 0;
        pixel_data[82][109] = 0;
        pixel_data[82][110] = 0;
        pixel_data[82][111] = 0;
        pixel_data[82][112] = 0;
        pixel_data[82][113] = 0;
        pixel_data[82][114] = 0;
        pixel_data[82][115] = 0;
        pixel_data[82][116] = 0;
        pixel_data[82][117] = 0;
        pixel_data[82][118] = 0;
        pixel_data[82][119] = 0;
        pixel_data[82][120] = 0;
        pixel_data[82][121] = 0;
        pixel_data[82][122] = 0;
        pixel_data[82][123] = 0;
        pixel_data[82][124] = 0;
        pixel_data[82][125] = 0;
        pixel_data[82][126] = 0;
        pixel_data[82][127] = 0;
        pixel_data[82][128] = 0;
        pixel_data[82][129] = 0;
        pixel_data[82][130] = 0;
        pixel_data[82][131] = 0;
        pixel_data[82][132] = 0;
        pixel_data[82][133] = 0;
        pixel_data[82][134] = 0;
        pixel_data[82][135] = 0;
        pixel_data[82][136] = 0;
        pixel_data[82][137] = 0;
        pixel_data[82][138] = 0;
        pixel_data[82][139] = 0;
        pixel_data[82][140] = 0;
        pixel_data[82][141] = 0;
        pixel_data[82][142] = 0;
        pixel_data[82][143] = 0;
        pixel_data[82][144] = 0;
        pixel_data[82][145] = 0;
        pixel_data[82][146] = 0;
        pixel_data[82][147] = 0;
        pixel_data[82][148] = 0;
        pixel_data[82][149] = 0;
        pixel_data[82][150] = 0;
        pixel_data[82][151] = 0;
        pixel_data[82][152] = 0;
        pixel_data[82][153] = 0;
        pixel_data[82][154] = 0;
        pixel_data[82][155] = 0;
        pixel_data[82][156] = 0;
        pixel_data[82][157] = 0;
        pixel_data[82][158] = 0;
        pixel_data[82][159] = 0;
        pixel_data[82][160] = 0;
        pixel_data[82][161] = 0;
        pixel_data[82][162] = 0;
        pixel_data[82][163] = 0;
        pixel_data[82][164] = 0;
        pixel_data[82][165] = 0;
        pixel_data[82][166] = 0;
        pixel_data[82][167] = 0;
        pixel_data[82][168] = 0;
        pixel_data[82][169] = 0;
        pixel_data[82][170] = 0;
        pixel_data[82][171] = 0;
        pixel_data[82][172] = 0;
        pixel_data[82][173] = 0;
        pixel_data[82][174] = 0;
        pixel_data[82][175] = 0;
        pixel_data[82][176] = 0;
        pixel_data[82][177] = 0;
        pixel_data[82][178] = 0;
        pixel_data[82][179] = 0;
        pixel_data[82][180] = 0;
        pixel_data[82][181] = 0;
        pixel_data[82][182] = 0;
        pixel_data[82][183] = 0;
        pixel_data[82][184] = 0;
        pixel_data[82][185] = 0;
        pixel_data[82][186] = 0;
        pixel_data[82][187] = 0;
        pixel_data[82][188] = 0;
        pixel_data[82][189] = 0;
        pixel_data[82][190] = 0;
        pixel_data[82][191] = 0;
        pixel_data[82][192] = 0;
        pixel_data[82][193] = 0;
        pixel_data[82][194] = 0;
        pixel_data[82][195] = 0;
        pixel_data[82][196] = 0;
        pixel_data[82][197] = 0;
        pixel_data[82][198] = 0;
        pixel_data[82][199] = 0; // y=82
        pixel_data[83][0] = 0;
        pixel_data[83][1] = 0;
        pixel_data[83][2] = 0;
        pixel_data[83][3] = 0;
        pixel_data[83][4] = 0;
        pixel_data[83][5] = 0;
        pixel_data[83][6] = 0;
        pixel_data[83][7] = 0;
        pixel_data[83][8] = 0;
        pixel_data[83][9] = 0;
        pixel_data[83][10] = 0;
        pixel_data[83][11] = 0;
        pixel_data[83][12] = 0;
        pixel_data[83][13] = 0;
        pixel_data[83][14] = 0;
        pixel_data[83][15] = 0;
        pixel_data[83][16] = 0;
        pixel_data[83][17] = 0;
        pixel_data[83][18] = 0;
        pixel_data[83][19] = 0;
        pixel_data[83][20] = 0;
        pixel_data[83][21] = 0;
        pixel_data[83][22] = 0;
        pixel_data[83][23] = 0;
        pixel_data[83][24] = 0;
        pixel_data[83][25] = 0;
        pixel_data[83][26] = 0;
        pixel_data[83][27] = 0;
        pixel_data[83][28] = 0;
        pixel_data[83][29] = 0;
        pixel_data[83][30] = 0;
        pixel_data[83][31] = 0;
        pixel_data[83][32] = 0;
        pixel_data[83][33] = 0;
        pixel_data[83][34] = 0;
        pixel_data[83][35] = 0;
        pixel_data[83][36] = 0;
        pixel_data[83][37] = 0;
        pixel_data[83][38] = 0;
        pixel_data[83][39] = 0;
        pixel_data[83][40] = 0;
        pixel_data[83][41] = 0;
        pixel_data[83][42] = 0;
        pixel_data[83][43] = 0;
        pixel_data[83][44] = 0;
        pixel_data[83][45] = 0;
        pixel_data[83][46] = 0;
        pixel_data[83][47] = 0;
        pixel_data[83][48] = 0;
        pixel_data[83][49] = 0;
        pixel_data[83][50] = 0;
        pixel_data[83][51] = 0;
        pixel_data[83][52] = 0;
        pixel_data[83][53] = 0;
        pixel_data[83][54] = 0;
        pixel_data[83][55] = 0;
        pixel_data[83][56] = 0;
        pixel_data[83][57] = 0;
        pixel_data[83][58] = 0;
        pixel_data[83][59] = 0;
        pixel_data[83][60] = 0;
        pixel_data[83][61] = 0;
        pixel_data[83][62] = 0;
        pixel_data[83][63] = 0;
        pixel_data[83][64] = 0;
        pixel_data[83][65] = 0;
        pixel_data[83][66] = 0;
        pixel_data[83][67] = 0;
        pixel_data[83][68] = 0;
        pixel_data[83][69] = 0;
        pixel_data[83][70] = 0;
        pixel_data[83][71] = 0;
        pixel_data[83][72] = 0;
        pixel_data[83][73] = 0;
        pixel_data[83][74] = 0;
        pixel_data[83][75] = 0;
        pixel_data[83][76] = 0;
        pixel_data[83][77] = 0;
        pixel_data[83][78] = 0;
        pixel_data[83][79] = 0;
        pixel_data[83][80] = 0;
        pixel_data[83][81] = 0;
        pixel_data[83][82] = 0;
        pixel_data[83][83] = 0;
        pixel_data[83][84] = 0;
        pixel_data[83][85] = 0;
        pixel_data[83][86] = 0;
        pixel_data[83][87] = 0;
        pixel_data[83][88] = 0;
        pixel_data[83][89] = 0;
        pixel_data[83][90] = 0;
        pixel_data[83][91] = 0;
        pixel_data[83][92] = 0;
        pixel_data[83][93] = 0;
        pixel_data[83][94] = 0;
        pixel_data[83][95] = 0;
        pixel_data[83][96] = 0;
        pixel_data[83][97] = 0;
        pixel_data[83][98] = 0;
        pixel_data[83][99] = 0;
        pixel_data[83][100] = 0;
        pixel_data[83][101] = 0;
        pixel_data[83][102] = 0;
        pixel_data[83][103] = 0;
        pixel_data[83][104] = 0;
        pixel_data[83][105] = 0;
        pixel_data[83][106] = 0;
        pixel_data[83][107] = 0;
        pixel_data[83][108] = 0;
        pixel_data[83][109] = 0;
        pixel_data[83][110] = 0;
        pixel_data[83][111] = 0;
        pixel_data[83][112] = 0;
        pixel_data[83][113] = 0;
        pixel_data[83][114] = 0;
        pixel_data[83][115] = 0;
        pixel_data[83][116] = 0;
        pixel_data[83][117] = 0;
        pixel_data[83][118] = 0;
        pixel_data[83][119] = 0;
        pixel_data[83][120] = 0;
        pixel_data[83][121] = 0;
        pixel_data[83][122] = 0;
        pixel_data[83][123] = 0;
        pixel_data[83][124] = 0;
        pixel_data[83][125] = 0;
        pixel_data[83][126] = 0;
        pixel_data[83][127] = 0;
        pixel_data[83][128] = 0;
        pixel_data[83][129] = 0;
        pixel_data[83][130] = 0;
        pixel_data[83][131] = 0;
        pixel_data[83][132] = 0;
        pixel_data[83][133] = 0;
        pixel_data[83][134] = 0;
        pixel_data[83][135] = 0;
        pixel_data[83][136] = 0;
        pixel_data[83][137] = 0;
        pixel_data[83][138] = 0;
        pixel_data[83][139] = 0;
        pixel_data[83][140] = 0;
        pixel_data[83][141] = 0;
        pixel_data[83][142] = 0;
        pixel_data[83][143] = 0;
        pixel_data[83][144] = 0;
        pixel_data[83][145] = 0;
        pixel_data[83][146] = 0;
        pixel_data[83][147] = 0;
        pixel_data[83][148] = 0;
        pixel_data[83][149] = 0;
        pixel_data[83][150] = 0;
        pixel_data[83][151] = 0;
        pixel_data[83][152] = 0;
        pixel_data[83][153] = 0;
        pixel_data[83][154] = 0;
        pixel_data[83][155] = 0;
        pixel_data[83][156] = 0;
        pixel_data[83][157] = 0;
        pixel_data[83][158] = 0;
        pixel_data[83][159] = 0;
        pixel_data[83][160] = 0;
        pixel_data[83][161] = 0;
        pixel_data[83][162] = 0;
        pixel_data[83][163] = 0;
        pixel_data[83][164] = 0;
        pixel_data[83][165] = 0;
        pixel_data[83][166] = 0;
        pixel_data[83][167] = 0;
        pixel_data[83][168] = 0;
        pixel_data[83][169] = 0;
        pixel_data[83][170] = 0;
        pixel_data[83][171] = 0;
        pixel_data[83][172] = 0;
        pixel_data[83][173] = 0;
        pixel_data[83][174] = 0;
        pixel_data[83][175] = 0;
        pixel_data[83][176] = 0;
        pixel_data[83][177] = 0;
        pixel_data[83][178] = 0;
        pixel_data[83][179] = 0;
        pixel_data[83][180] = 0;
        pixel_data[83][181] = 0;
        pixel_data[83][182] = 0;
        pixel_data[83][183] = 0;
        pixel_data[83][184] = 0;
        pixel_data[83][185] = 0;
        pixel_data[83][186] = 0;
        pixel_data[83][187] = 0;
        pixel_data[83][188] = 0;
        pixel_data[83][189] = 0;
        pixel_data[83][190] = 0;
        pixel_data[83][191] = 0;
        pixel_data[83][192] = 0;
        pixel_data[83][193] = 0;
        pixel_data[83][194] = 0;
        pixel_data[83][195] = 0;
        pixel_data[83][196] = 0;
        pixel_data[83][197] = 0;
        pixel_data[83][198] = 0;
        pixel_data[83][199] = 0; // y=83
        pixel_data[84][0] = 0;
        pixel_data[84][1] = 0;
        pixel_data[84][2] = 0;
        pixel_data[84][3] = 0;
        pixel_data[84][4] = 0;
        pixel_data[84][5] = 0;
        pixel_data[84][6] = 0;
        pixel_data[84][7] = 0;
        pixel_data[84][8] = 0;
        pixel_data[84][9] = 0;
        pixel_data[84][10] = 0;
        pixel_data[84][11] = 0;
        pixel_data[84][12] = 0;
        pixel_data[84][13] = 0;
        pixel_data[84][14] = 0;
        pixel_data[84][15] = 0;
        pixel_data[84][16] = 0;
        pixel_data[84][17] = 0;
        pixel_data[84][18] = 0;
        pixel_data[84][19] = 0;
        pixel_data[84][20] = 0;
        pixel_data[84][21] = 0;
        pixel_data[84][22] = 0;
        pixel_data[84][23] = 0;
        pixel_data[84][24] = 0;
        pixel_data[84][25] = 0;
        pixel_data[84][26] = 0;
        pixel_data[84][27] = 0;
        pixel_data[84][28] = 0;
        pixel_data[84][29] = 0;
        pixel_data[84][30] = 0;
        pixel_data[84][31] = 0;
        pixel_data[84][32] = 0;
        pixel_data[84][33] = 0;
        pixel_data[84][34] = 0;
        pixel_data[84][35] = 0;
        pixel_data[84][36] = 0;
        pixel_data[84][37] = 0;
        pixel_data[84][38] = 0;
        pixel_data[84][39] = 0;
        pixel_data[84][40] = 0;
        pixel_data[84][41] = 0;
        pixel_data[84][42] = 0;
        pixel_data[84][43] = 0;
        pixel_data[84][44] = 0;
        pixel_data[84][45] = 0;
        pixel_data[84][46] = 0;
        pixel_data[84][47] = 0;
        pixel_data[84][48] = 0;
        pixel_data[84][49] = 0;
        pixel_data[84][50] = 0;
        pixel_data[84][51] = 0;
        pixel_data[84][52] = 0;
        pixel_data[84][53] = 0;
        pixel_data[84][54] = 0;
        pixel_data[84][55] = 0;
        pixel_data[84][56] = 0;
        pixel_data[84][57] = 0;
        pixel_data[84][58] = 0;
        pixel_data[84][59] = 0;
        pixel_data[84][60] = 0;
        pixel_data[84][61] = 0;
        pixel_data[84][62] = 0;
        pixel_data[84][63] = 0;
        pixel_data[84][64] = 0;
        pixel_data[84][65] = 0;
        pixel_data[84][66] = 0;
        pixel_data[84][67] = 0;
        pixel_data[84][68] = 0;
        pixel_data[84][69] = 0;
        pixel_data[84][70] = 0;
        pixel_data[84][71] = 0;
        pixel_data[84][72] = 0;
        pixel_data[84][73] = 0;
        pixel_data[84][74] = 0;
        pixel_data[84][75] = 0;
        pixel_data[84][76] = 0;
        pixel_data[84][77] = 0;
        pixel_data[84][78] = 0;
        pixel_data[84][79] = 0;
        pixel_data[84][80] = 0;
        pixel_data[84][81] = 0;
        pixel_data[84][82] = 0;
        pixel_data[84][83] = 0;
        pixel_data[84][84] = 0;
        pixel_data[84][85] = 0;
        pixel_data[84][86] = 0;
        pixel_data[84][87] = 0;
        pixel_data[84][88] = 0;
        pixel_data[84][89] = 0;
        pixel_data[84][90] = 0;
        pixel_data[84][91] = 0;
        pixel_data[84][92] = 0;
        pixel_data[84][93] = 0;
        pixel_data[84][94] = 0;
        pixel_data[84][95] = 0;
        pixel_data[84][96] = 0;
        pixel_data[84][97] = 0;
        pixel_data[84][98] = 0;
        pixel_data[84][99] = 0;
        pixel_data[84][100] = 0;
        pixel_data[84][101] = 0;
        pixel_data[84][102] = 0;
        pixel_data[84][103] = 0;
        pixel_data[84][104] = 0;
        pixel_data[84][105] = 0;
        pixel_data[84][106] = 0;
        pixel_data[84][107] = 0;
        pixel_data[84][108] = 0;
        pixel_data[84][109] = 0;
        pixel_data[84][110] = 0;
        pixel_data[84][111] = 0;
        pixel_data[84][112] = 0;
        pixel_data[84][113] = 0;
        pixel_data[84][114] = 0;
        pixel_data[84][115] = 0;
        pixel_data[84][116] = 0;
        pixel_data[84][117] = 0;
        pixel_data[84][118] = 0;
        pixel_data[84][119] = 0;
        pixel_data[84][120] = 0;
        pixel_data[84][121] = 0;
        pixel_data[84][122] = 0;
        pixel_data[84][123] = 0;
        pixel_data[84][124] = 0;
        pixel_data[84][125] = 0;
        pixel_data[84][126] = 0;
        pixel_data[84][127] = 0;
        pixel_data[84][128] = 0;
        pixel_data[84][129] = 0;
        pixel_data[84][130] = 0;
        pixel_data[84][131] = 0;
        pixel_data[84][132] = 0;
        pixel_data[84][133] = 0;
        pixel_data[84][134] = 0;
        pixel_data[84][135] = 0;
        pixel_data[84][136] = 0;
        pixel_data[84][137] = 0;
        pixel_data[84][138] = 0;
        pixel_data[84][139] = 0;
        pixel_data[84][140] = 0;
        pixel_data[84][141] = 0;
        pixel_data[84][142] = 0;
        pixel_data[84][143] = 0;
        pixel_data[84][144] = 0;
        pixel_data[84][145] = 0;
        pixel_data[84][146] = 0;
        pixel_data[84][147] = 0;
        pixel_data[84][148] = 0;
        pixel_data[84][149] = 0;
        pixel_data[84][150] = 0;
        pixel_data[84][151] = 0;
        pixel_data[84][152] = 0;
        pixel_data[84][153] = 0;
        pixel_data[84][154] = 0;
        pixel_data[84][155] = 0;
        pixel_data[84][156] = 0;
        pixel_data[84][157] = 0;
        pixel_data[84][158] = 0;
        pixel_data[84][159] = 0;
        pixel_data[84][160] = 0;
        pixel_data[84][161] = 0;
        pixel_data[84][162] = 0;
        pixel_data[84][163] = 0;
        pixel_data[84][164] = 0;
        pixel_data[84][165] = 0;
        pixel_data[84][166] = 0;
        pixel_data[84][167] = 0;
        pixel_data[84][168] = 0;
        pixel_data[84][169] = 0;
        pixel_data[84][170] = 0;
        pixel_data[84][171] = 0;
        pixel_data[84][172] = 0;
        pixel_data[84][173] = 0;
        pixel_data[84][174] = 0;
        pixel_data[84][175] = 0;
        pixel_data[84][176] = 0;
        pixel_data[84][177] = 0;
        pixel_data[84][178] = 0;
        pixel_data[84][179] = 0;
        pixel_data[84][180] = 0;
        pixel_data[84][181] = 0;
        pixel_data[84][182] = 0;
        pixel_data[84][183] = 0;
        pixel_data[84][184] = 0;
        pixel_data[84][185] = 0;
        pixel_data[84][186] = 0;
        pixel_data[84][187] = 0;
        pixel_data[84][188] = 0;
        pixel_data[84][189] = 0;
        pixel_data[84][190] = 0;
        pixel_data[84][191] = 0;
        pixel_data[84][192] = 0;
        pixel_data[84][193] = 0;
        pixel_data[84][194] = 0;
        pixel_data[84][195] = 0;
        pixel_data[84][196] = 0;
        pixel_data[84][197] = 0;
        pixel_data[84][198] = 0;
        pixel_data[84][199] = 0; // y=84
        pixel_data[85][0] = 0;
        pixel_data[85][1] = 0;
        pixel_data[85][2] = 0;
        pixel_data[85][3] = 0;
        pixel_data[85][4] = 0;
        pixel_data[85][5] = 0;
        pixel_data[85][6] = 0;
        pixel_data[85][7] = 0;
        pixel_data[85][8] = 0;
        pixel_data[85][9] = 0;
        pixel_data[85][10] = 0;
        pixel_data[85][11] = 0;
        pixel_data[85][12] = 0;
        pixel_data[85][13] = 0;
        pixel_data[85][14] = 0;
        pixel_data[85][15] = 0;
        pixel_data[85][16] = 0;
        pixel_data[85][17] = 0;
        pixel_data[85][18] = 0;
        pixel_data[85][19] = 0;
        pixel_data[85][20] = 0;
        pixel_data[85][21] = 0;
        pixel_data[85][22] = 0;
        pixel_data[85][23] = 0;
        pixel_data[85][24] = 0;
        pixel_data[85][25] = 0;
        pixel_data[85][26] = 0;
        pixel_data[85][27] = 0;
        pixel_data[85][28] = 0;
        pixel_data[85][29] = 0;
        pixel_data[85][30] = 0;
        pixel_data[85][31] = 0;
        pixel_data[85][32] = 0;
        pixel_data[85][33] = 0;
        pixel_data[85][34] = 0;
        pixel_data[85][35] = 0;
        pixel_data[85][36] = 0;
        pixel_data[85][37] = 0;
        pixel_data[85][38] = 0;
        pixel_data[85][39] = 0;
        pixel_data[85][40] = 0;
        pixel_data[85][41] = 0;
        pixel_data[85][42] = 0;
        pixel_data[85][43] = 0;
        pixel_data[85][44] = 0;
        pixel_data[85][45] = 0;
        pixel_data[85][46] = 0;
        pixel_data[85][47] = 0;
        pixel_data[85][48] = 0;
        pixel_data[85][49] = 0;
        pixel_data[85][50] = 0;
        pixel_data[85][51] = 0;
        pixel_data[85][52] = 0;
        pixel_data[85][53] = 0;
        pixel_data[85][54] = 0;
        pixel_data[85][55] = 0;
        pixel_data[85][56] = 0;
        pixel_data[85][57] = 0;
        pixel_data[85][58] = 0;
        pixel_data[85][59] = 0;
        pixel_data[85][60] = 0;
        pixel_data[85][61] = 0;
        pixel_data[85][62] = 0;
        pixel_data[85][63] = 0;
        pixel_data[85][64] = 0;
        pixel_data[85][65] = 0;
        pixel_data[85][66] = 0;
        pixel_data[85][67] = 0;
        pixel_data[85][68] = 0;
        pixel_data[85][69] = 0;
        pixel_data[85][70] = 0;
        pixel_data[85][71] = 0;
        pixel_data[85][72] = 0;
        pixel_data[85][73] = 0;
        pixel_data[85][74] = 0;
        pixel_data[85][75] = 0;
        pixel_data[85][76] = 0;
        pixel_data[85][77] = 0;
        pixel_data[85][78] = 0;
        pixel_data[85][79] = 0;
        pixel_data[85][80] = 0;
        pixel_data[85][81] = 0;
        pixel_data[85][82] = 0;
        pixel_data[85][83] = 0;
        pixel_data[85][84] = 0;
        pixel_data[85][85] = 0;
        pixel_data[85][86] = 0;
        pixel_data[85][87] = 0;
        pixel_data[85][88] = 0;
        pixel_data[85][89] = 0;
        pixel_data[85][90] = 0;
        pixel_data[85][91] = 0;
        pixel_data[85][92] = 0;
        pixel_data[85][93] = 0;
        pixel_data[85][94] = 0;
        pixel_data[85][95] = 0;
        pixel_data[85][96] = 0;
        pixel_data[85][97] = 0;
        pixel_data[85][98] = 0;
        pixel_data[85][99] = 0;
        pixel_data[85][100] = 0;
        pixel_data[85][101] = 0;
        pixel_data[85][102] = 0;
        pixel_data[85][103] = 0;
        pixel_data[85][104] = 0;
        pixel_data[85][105] = 0;
        pixel_data[85][106] = 0;
        pixel_data[85][107] = 0;
        pixel_data[85][108] = 0;
        pixel_data[85][109] = 0;
        pixel_data[85][110] = 0;
        pixel_data[85][111] = 0;
        pixel_data[85][112] = 0;
        pixel_data[85][113] = 0;
        pixel_data[85][114] = 0;
        pixel_data[85][115] = 0;
        pixel_data[85][116] = 0;
        pixel_data[85][117] = 0;
        pixel_data[85][118] = 0;
        pixel_data[85][119] = 0;
        pixel_data[85][120] = 0;
        pixel_data[85][121] = 0;
        pixel_data[85][122] = 0;
        pixel_data[85][123] = 0;
        pixel_data[85][124] = 0;
        pixel_data[85][125] = 0;
        pixel_data[85][126] = 0;
        pixel_data[85][127] = 0;
        pixel_data[85][128] = 0;
        pixel_data[85][129] = 0;
        pixel_data[85][130] = 0;
        pixel_data[85][131] = 0;
        pixel_data[85][132] = 0;
        pixel_data[85][133] = 0;
        pixel_data[85][134] = 0;
        pixel_data[85][135] = 0;
        pixel_data[85][136] = 0;
        pixel_data[85][137] = 0;
        pixel_data[85][138] = 0;
        pixel_data[85][139] = 0;
        pixel_data[85][140] = 0;
        pixel_data[85][141] = 0;
        pixel_data[85][142] = 0;
        pixel_data[85][143] = 0;
        pixel_data[85][144] = 0;
        pixel_data[85][145] = 0;
        pixel_data[85][146] = 0;
        pixel_data[85][147] = 0;
        pixel_data[85][148] = 0;
        pixel_data[85][149] = 0;
        pixel_data[85][150] = 0;
        pixel_data[85][151] = 0;
        pixel_data[85][152] = 0;
        pixel_data[85][153] = 0;
        pixel_data[85][154] = 0;
        pixel_data[85][155] = 0;
        pixel_data[85][156] = 0;
        pixel_data[85][157] = 0;
        pixel_data[85][158] = 0;
        pixel_data[85][159] = 0;
        pixel_data[85][160] = 0;
        pixel_data[85][161] = 0;
        pixel_data[85][162] = 0;
        pixel_data[85][163] = 0;
        pixel_data[85][164] = 0;
        pixel_data[85][165] = 0;
        pixel_data[85][166] = 0;
        pixel_data[85][167] = 0;
        pixel_data[85][168] = 0;
        pixel_data[85][169] = 0;
        pixel_data[85][170] = 0;
        pixel_data[85][171] = 0;
        pixel_data[85][172] = 0;
        pixel_data[85][173] = 0;
        pixel_data[85][174] = 0;
        pixel_data[85][175] = 0;
        pixel_data[85][176] = 0;
        pixel_data[85][177] = 0;
        pixel_data[85][178] = 0;
        pixel_data[85][179] = 0;
        pixel_data[85][180] = 0;
        pixel_data[85][181] = 0;
        pixel_data[85][182] = 0;
        pixel_data[85][183] = 0;
        pixel_data[85][184] = 0;
        pixel_data[85][185] = 0;
        pixel_data[85][186] = 0;
        pixel_data[85][187] = 0;
        pixel_data[85][188] = 0;
        pixel_data[85][189] = 0;
        pixel_data[85][190] = 0;
        pixel_data[85][191] = 0;
        pixel_data[85][192] = 0;
        pixel_data[85][193] = 0;
        pixel_data[85][194] = 0;
        pixel_data[85][195] = 0;
        pixel_data[85][196] = 0;
        pixel_data[85][197] = 0;
        pixel_data[85][198] = 0;
        pixel_data[85][199] = 0; // y=85
        pixel_data[86][0] = 0;
        pixel_data[86][1] = 0;
        pixel_data[86][2] = 0;
        pixel_data[86][3] = 0;
        pixel_data[86][4] = 0;
        pixel_data[86][5] = 0;
        pixel_data[86][6] = 0;
        pixel_data[86][7] = 0;
        pixel_data[86][8] = 0;
        pixel_data[86][9] = 0;
        pixel_data[86][10] = 0;
        pixel_data[86][11] = 0;
        pixel_data[86][12] = 0;
        pixel_data[86][13] = 0;
        pixel_data[86][14] = 0;
        pixel_data[86][15] = 0;
        pixel_data[86][16] = 0;
        pixel_data[86][17] = 0;
        pixel_data[86][18] = 0;
        pixel_data[86][19] = 0;
        pixel_data[86][20] = 0;
        pixel_data[86][21] = 0;
        pixel_data[86][22] = 0;
        pixel_data[86][23] = 0;
        pixel_data[86][24] = 0;
        pixel_data[86][25] = 0;
        pixel_data[86][26] = 0;
        pixel_data[86][27] = 0;
        pixel_data[86][28] = 0;
        pixel_data[86][29] = 0;
        pixel_data[86][30] = 0;
        pixel_data[86][31] = 0;
        pixel_data[86][32] = 0;
        pixel_data[86][33] = 0;
        pixel_data[86][34] = 0;
        pixel_data[86][35] = 0;
        pixel_data[86][36] = 0;
        pixel_data[86][37] = 0;
        pixel_data[86][38] = 0;
        pixel_data[86][39] = 0;
        pixel_data[86][40] = 0;
        pixel_data[86][41] = 0;
        pixel_data[86][42] = 0;
        pixel_data[86][43] = 0;
        pixel_data[86][44] = 0;
        pixel_data[86][45] = 0;
        pixel_data[86][46] = 0;
        pixel_data[86][47] = 0;
        pixel_data[86][48] = 0;
        pixel_data[86][49] = 0;
        pixel_data[86][50] = 0;
        pixel_data[86][51] = 0;
        pixel_data[86][52] = 0;
        pixel_data[86][53] = 0;
        pixel_data[86][54] = 0;
        pixel_data[86][55] = 0;
        pixel_data[86][56] = 0;
        pixel_data[86][57] = 0;
        pixel_data[86][58] = 0;
        pixel_data[86][59] = 0;
        pixel_data[86][60] = 0;
        pixel_data[86][61] = 0;
        pixel_data[86][62] = 0;
        pixel_data[86][63] = 0;
        pixel_data[86][64] = 0;
        pixel_data[86][65] = 0;
        pixel_data[86][66] = 0;
        pixel_data[86][67] = 0;
        pixel_data[86][68] = 0;
        pixel_data[86][69] = 0;
        pixel_data[86][70] = 0;
        pixel_data[86][71] = 0;
        pixel_data[86][72] = 0;
        pixel_data[86][73] = 0;
        pixel_data[86][74] = 0;
        pixel_data[86][75] = 0;
        pixel_data[86][76] = 0;
        pixel_data[86][77] = 0;
        pixel_data[86][78] = 0;
        pixel_data[86][79] = 0;
        pixel_data[86][80] = 0;
        pixel_data[86][81] = 0;
        pixel_data[86][82] = 0;
        pixel_data[86][83] = 0;
        pixel_data[86][84] = 0;
        pixel_data[86][85] = 0;
        pixel_data[86][86] = 0;
        pixel_data[86][87] = 0;
        pixel_data[86][88] = 0;
        pixel_data[86][89] = 0;
        pixel_data[86][90] = 0;
        pixel_data[86][91] = 0;
        pixel_data[86][92] = 0;
        pixel_data[86][93] = 0;
        pixel_data[86][94] = 0;
        pixel_data[86][95] = 0;
        pixel_data[86][96] = 0;
        pixel_data[86][97] = 0;
        pixel_data[86][98] = 0;
        pixel_data[86][99] = 0;
        pixel_data[86][100] = 0;
        pixel_data[86][101] = 0;
        pixel_data[86][102] = 0;
        pixel_data[86][103] = 0;
        pixel_data[86][104] = 0;
        pixel_data[86][105] = 0;
        pixel_data[86][106] = 0;
        pixel_data[86][107] = 0;
        pixel_data[86][108] = 0;
        pixel_data[86][109] = 0;
        pixel_data[86][110] = 0;
        pixel_data[86][111] = 0;
        pixel_data[86][112] = 0;
        pixel_data[86][113] = 0;
        pixel_data[86][114] = 0;
        pixel_data[86][115] = 0;
        pixel_data[86][116] = 0;
        pixel_data[86][117] = 0;
        pixel_data[86][118] = 0;
        pixel_data[86][119] = 0;
        pixel_data[86][120] = 0;
        pixel_data[86][121] = 0;
        pixel_data[86][122] = 0;
        pixel_data[86][123] = 0;
        pixel_data[86][124] = 0;
        pixel_data[86][125] = 0;
        pixel_data[86][126] = 0;
        pixel_data[86][127] = 0;
        pixel_data[86][128] = 0;
        pixel_data[86][129] = 0;
        pixel_data[86][130] = 0;
        pixel_data[86][131] = 0;
        pixel_data[86][132] = 0;
        pixel_data[86][133] = 0;
        pixel_data[86][134] = 0;
        pixel_data[86][135] = 0;
        pixel_data[86][136] = 0;
        pixel_data[86][137] = 0;
        pixel_data[86][138] = 0;
        pixel_data[86][139] = 0;
        pixel_data[86][140] = 0;
        pixel_data[86][141] = 0;
        pixel_data[86][142] = 0;
        pixel_data[86][143] = 0;
        pixel_data[86][144] = 0;
        pixel_data[86][145] = 0;
        pixel_data[86][146] = 0;
        pixel_data[86][147] = 0;
        pixel_data[86][148] = 0;
        pixel_data[86][149] = 0;
        pixel_data[86][150] = 0;
        pixel_data[86][151] = 0;
        pixel_data[86][152] = 0;
        pixel_data[86][153] = 0;
        pixel_data[86][154] = 0;
        pixel_data[86][155] = 0;
        pixel_data[86][156] = 0;
        pixel_data[86][157] = 0;
        pixel_data[86][158] = 0;
        pixel_data[86][159] = 0;
        pixel_data[86][160] = 0;
        pixel_data[86][161] = 0;
        pixel_data[86][162] = 0;
        pixel_data[86][163] = 0;
        pixel_data[86][164] = 0;
        pixel_data[86][165] = 0;
        pixel_data[86][166] = 0;
        pixel_data[86][167] = 0;
        pixel_data[86][168] = 0;
        pixel_data[86][169] = 0;
        pixel_data[86][170] = 0;
        pixel_data[86][171] = 0;
        pixel_data[86][172] = 0;
        pixel_data[86][173] = 0;
        pixel_data[86][174] = 0;
        pixel_data[86][175] = 0;
        pixel_data[86][176] = 0;
        pixel_data[86][177] = 0;
        pixel_data[86][178] = 0;
        pixel_data[86][179] = 0;
        pixel_data[86][180] = 0;
        pixel_data[86][181] = 0;
        pixel_data[86][182] = 0;
        pixel_data[86][183] = 0;
        pixel_data[86][184] = 0;
        pixel_data[86][185] = 0;
        pixel_data[86][186] = 0;
        pixel_data[86][187] = 0;
        pixel_data[86][188] = 0;
        pixel_data[86][189] = 0;
        pixel_data[86][190] = 0;
        pixel_data[86][191] = 0;
        pixel_data[86][192] = 0;
        pixel_data[86][193] = 0;
        pixel_data[86][194] = 0;
        pixel_data[86][195] = 0;
        pixel_data[86][196] = 0;
        pixel_data[86][197] = 0;
        pixel_data[86][198] = 0;
        pixel_data[86][199] = 0; // y=86
        pixel_data[87][0] = 0;
        pixel_data[87][1] = 0;
        pixel_data[87][2] = 0;
        pixel_data[87][3] = 0;
        pixel_data[87][4] = 0;
        pixel_data[87][5] = 0;
        pixel_data[87][6] = 0;
        pixel_data[87][7] = 0;
        pixel_data[87][8] = 0;
        pixel_data[87][9] = 0;
        pixel_data[87][10] = 0;
        pixel_data[87][11] = 0;
        pixel_data[87][12] = 0;
        pixel_data[87][13] = 0;
        pixel_data[87][14] = 0;
        pixel_data[87][15] = 0;
        pixel_data[87][16] = 0;
        pixel_data[87][17] = 0;
        pixel_data[87][18] = 0;
        pixel_data[87][19] = 0;
        pixel_data[87][20] = 0;
        pixel_data[87][21] = 0;
        pixel_data[87][22] = 0;
        pixel_data[87][23] = 0;
        pixel_data[87][24] = 0;
        pixel_data[87][25] = 0;
        pixel_data[87][26] = 0;
        pixel_data[87][27] = 0;
        pixel_data[87][28] = 0;
        pixel_data[87][29] = 0;
        pixel_data[87][30] = 0;
        pixel_data[87][31] = 0;
        pixel_data[87][32] = 0;
        pixel_data[87][33] = 0;
        pixel_data[87][34] = 0;
        pixel_data[87][35] = 0;
        pixel_data[87][36] = 0;
        pixel_data[87][37] = 0;
        pixel_data[87][38] = 0;
        pixel_data[87][39] = 0;
        pixel_data[87][40] = 0;
        pixel_data[87][41] = 0;
        pixel_data[87][42] = 0;
        pixel_data[87][43] = 0;
        pixel_data[87][44] = 0;
        pixel_data[87][45] = 0;
        pixel_data[87][46] = 0;
        pixel_data[87][47] = 0;
        pixel_data[87][48] = 0;
        pixel_data[87][49] = 0;
        pixel_data[87][50] = 0;
        pixel_data[87][51] = 0;
        pixel_data[87][52] = 0;
        pixel_data[87][53] = 0;
        pixel_data[87][54] = 0;
        pixel_data[87][55] = 0;
        pixel_data[87][56] = 0;
        pixel_data[87][57] = 0;
        pixel_data[87][58] = 0;
        pixel_data[87][59] = 0;
        pixel_data[87][60] = 0;
        pixel_data[87][61] = 0;
        pixel_data[87][62] = 0;
        pixel_data[87][63] = 0;
        pixel_data[87][64] = 0;
        pixel_data[87][65] = 0;
        pixel_data[87][66] = 0;
        pixel_data[87][67] = 0;
        pixel_data[87][68] = 0;
        pixel_data[87][69] = 0;
        pixel_data[87][70] = 0;
        pixel_data[87][71] = 0;
        pixel_data[87][72] = 0;
        pixel_data[87][73] = 0;
        pixel_data[87][74] = 0;
        pixel_data[87][75] = 0;
        pixel_data[87][76] = 0;
        pixel_data[87][77] = 0;
        pixel_data[87][78] = 0;
        pixel_data[87][79] = 0;
        pixel_data[87][80] = 0;
        pixel_data[87][81] = 0;
        pixel_data[87][82] = 0;
        pixel_data[87][83] = 0;
        pixel_data[87][84] = 0;
        pixel_data[87][85] = 0;
        pixel_data[87][86] = 0;
        pixel_data[87][87] = 0;
        pixel_data[87][88] = 0;
        pixel_data[87][89] = 0;
        pixel_data[87][90] = 0;
        pixel_data[87][91] = 0;
        pixel_data[87][92] = 0;
        pixel_data[87][93] = 0;
        pixel_data[87][94] = 0;
        pixel_data[87][95] = 0;
        pixel_data[87][96] = 0;
        pixel_data[87][97] = 0;
        pixel_data[87][98] = 0;
        pixel_data[87][99] = 0;
        pixel_data[87][100] = 0;
        pixel_data[87][101] = 0;
        pixel_data[87][102] = 0;
        pixel_data[87][103] = 0;
        pixel_data[87][104] = 0;
        pixel_data[87][105] = 0;
        pixel_data[87][106] = 0;
        pixel_data[87][107] = 0;
        pixel_data[87][108] = 0;
        pixel_data[87][109] = 0;
        pixel_data[87][110] = 0;
        pixel_data[87][111] = 0;
        pixel_data[87][112] = 0;
        pixel_data[87][113] = 0;
        pixel_data[87][114] = 0;
        pixel_data[87][115] = 0;
        pixel_data[87][116] = 0;
        pixel_data[87][117] = 0;
        pixel_data[87][118] = 0;
        pixel_data[87][119] = 0;
        pixel_data[87][120] = 0;
        pixel_data[87][121] = 0;
        pixel_data[87][122] = 0;
        pixel_data[87][123] = 0;
        pixel_data[87][124] = 0;
        pixel_data[87][125] = 0;
        pixel_data[87][126] = 0;
        pixel_data[87][127] = 0;
        pixel_data[87][128] = 0;
        pixel_data[87][129] = 0;
        pixel_data[87][130] = 0;
        pixel_data[87][131] = 0;
        pixel_data[87][132] = 0;
        pixel_data[87][133] = 0;
        pixel_data[87][134] = 0;
        pixel_data[87][135] = 0;
        pixel_data[87][136] = 0;
        pixel_data[87][137] = 0;
        pixel_data[87][138] = 0;
        pixel_data[87][139] = 0;
        pixel_data[87][140] = 0;
        pixel_data[87][141] = 0;
        pixel_data[87][142] = 0;
        pixel_data[87][143] = 0;
        pixel_data[87][144] = 0;
        pixel_data[87][145] = 0;
        pixel_data[87][146] = 0;
        pixel_data[87][147] = 0;
        pixel_data[87][148] = 0;
        pixel_data[87][149] = 0;
        pixel_data[87][150] = 0;
        pixel_data[87][151] = 0;
        pixel_data[87][152] = 0;
        pixel_data[87][153] = 0;
        pixel_data[87][154] = 0;
        pixel_data[87][155] = 0;
        pixel_data[87][156] = 0;
        pixel_data[87][157] = 0;
        pixel_data[87][158] = 0;
        pixel_data[87][159] = 0;
        pixel_data[87][160] = 0;
        pixel_data[87][161] = 0;
        pixel_data[87][162] = 0;
        pixel_data[87][163] = 0;
        pixel_data[87][164] = 0;
        pixel_data[87][165] = 0;
        pixel_data[87][166] = 0;
        pixel_data[87][167] = 0;
        pixel_data[87][168] = 0;
        pixel_data[87][169] = 0;
        pixel_data[87][170] = 0;
        pixel_data[87][171] = 0;
        pixel_data[87][172] = 0;
        pixel_data[87][173] = 0;
        pixel_data[87][174] = 0;
        pixel_data[87][175] = 0;
        pixel_data[87][176] = 0;
        pixel_data[87][177] = 0;
        pixel_data[87][178] = 0;
        pixel_data[87][179] = 0;
        pixel_data[87][180] = 0;
        pixel_data[87][181] = 0;
        pixel_data[87][182] = 0;
        pixel_data[87][183] = 0;
        pixel_data[87][184] = 0;
        pixel_data[87][185] = 0;
        pixel_data[87][186] = 0;
        pixel_data[87][187] = 0;
        pixel_data[87][188] = 0;
        pixel_data[87][189] = 0;
        pixel_data[87][190] = 0;
        pixel_data[87][191] = 0;
        pixel_data[87][192] = 0;
        pixel_data[87][193] = 0;
        pixel_data[87][194] = 0;
        pixel_data[87][195] = 0;
        pixel_data[87][196] = 0;
        pixel_data[87][197] = 0;
        pixel_data[87][198] = 0;
        pixel_data[87][199] = 0; // y=87
        pixel_data[88][0] = 0;
        pixel_data[88][1] = 0;
        pixel_data[88][2] = 0;
        pixel_data[88][3] = 0;
        pixel_data[88][4] = 0;
        pixel_data[88][5] = 0;
        pixel_data[88][6] = 0;
        pixel_data[88][7] = 0;
        pixel_data[88][8] = 0;
        pixel_data[88][9] = 0;
        pixel_data[88][10] = 0;
        pixel_data[88][11] = 0;
        pixel_data[88][12] = 0;
        pixel_data[88][13] = 0;
        pixel_data[88][14] = 0;
        pixel_data[88][15] = 0;
        pixel_data[88][16] = 0;
        pixel_data[88][17] = 0;
        pixel_data[88][18] = 0;
        pixel_data[88][19] = 0;
        pixel_data[88][20] = 0;
        pixel_data[88][21] = 0;
        pixel_data[88][22] = 0;
        pixel_data[88][23] = 0;
        pixel_data[88][24] = 0;
        pixel_data[88][25] = 0;
        pixel_data[88][26] = 0;
        pixel_data[88][27] = 0;
        pixel_data[88][28] = 0;
        pixel_data[88][29] = 0;
        pixel_data[88][30] = 0;
        pixel_data[88][31] = 0;
        pixel_data[88][32] = 0;
        pixel_data[88][33] = 0;
        pixel_data[88][34] = 0;
        pixel_data[88][35] = 0;
        pixel_data[88][36] = 0;
        pixel_data[88][37] = 0;
        pixel_data[88][38] = 0;
        pixel_data[88][39] = 0;
        pixel_data[88][40] = 0;
        pixel_data[88][41] = 0;
        pixel_data[88][42] = 0;
        pixel_data[88][43] = 0;
        pixel_data[88][44] = 0;
        pixel_data[88][45] = 0;
        pixel_data[88][46] = 0;
        pixel_data[88][47] = 0;
        pixel_data[88][48] = 0;
        pixel_data[88][49] = 0;
        pixel_data[88][50] = 0;
        pixel_data[88][51] = 0;
        pixel_data[88][52] = 0;
        pixel_data[88][53] = 0;
        pixel_data[88][54] = 0;
        pixel_data[88][55] = 0;
        pixel_data[88][56] = 0;
        pixel_data[88][57] = 0;
        pixel_data[88][58] = 0;
        pixel_data[88][59] = 0;
        pixel_data[88][60] = 0;
        pixel_data[88][61] = 0;
        pixel_data[88][62] = 0;
        pixel_data[88][63] = 0;
        pixel_data[88][64] = 0;
        pixel_data[88][65] = 0;
        pixel_data[88][66] = 0;
        pixel_data[88][67] = 0;
        pixel_data[88][68] = 0;
        pixel_data[88][69] = 0;
        pixel_data[88][70] = 0;
        pixel_data[88][71] = 0;
        pixel_data[88][72] = 0;
        pixel_data[88][73] = 0;
        pixel_data[88][74] = 0;
        pixel_data[88][75] = 0;
        pixel_data[88][76] = 0;
        pixel_data[88][77] = 0;
        pixel_data[88][78] = 0;
        pixel_data[88][79] = 0;
        pixel_data[88][80] = 0;
        pixel_data[88][81] = 0;
        pixel_data[88][82] = 0;
        pixel_data[88][83] = 0;
        pixel_data[88][84] = 0;
        pixel_data[88][85] = 0;
        pixel_data[88][86] = 0;
        pixel_data[88][87] = 0;
        pixel_data[88][88] = 0;
        pixel_data[88][89] = 0;
        pixel_data[88][90] = 0;
        pixel_data[88][91] = 0;
        pixel_data[88][92] = 0;
        pixel_data[88][93] = 0;
        pixel_data[88][94] = 0;
        pixel_data[88][95] = 0;
        pixel_data[88][96] = 0;
        pixel_data[88][97] = 0;
        pixel_data[88][98] = 0;
        pixel_data[88][99] = 0;
        pixel_data[88][100] = 0;
        pixel_data[88][101] = 0;
        pixel_data[88][102] = 0;
        pixel_data[88][103] = 0;
        pixel_data[88][104] = 0;
        pixel_data[88][105] = 0;
        pixel_data[88][106] = 0;
        pixel_data[88][107] = 0;
        pixel_data[88][108] = 0;
        pixel_data[88][109] = 0;
        pixel_data[88][110] = 0;
        pixel_data[88][111] = 0;
        pixel_data[88][112] = 0;
        pixel_data[88][113] = 0;
        pixel_data[88][114] = 0;
        pixel_data[88][115] = 0;
        pixel_data[88][116] = 0;
        pixel_data[88][117] = 0;
        pixel_data[88][118] = 0;
        pixel_data[88][119] = 0;
        pixel_data[88][120] = 0;
        pixel_data[88][121] = 0;
        pixel_data[88][122] = 0;
        pixel_data[88][123] = 0;
        pixel_data[88][124] = 0;
        pixel_data[88][125] = 0;
        pixel_data[88][126] = 0;
        pixel_data[88][127] = 0;
        pixel_data[88][128] = 0;
        pixel_data[88][129] = 0;
        pixel_data[88][130] = 0;
        pixel_data[88][131] = 0;
        pixel_data[88][132] = 0;
        pixel_data[88][133] = 0;
        pixel_data[88][134] = 0;
        pixel_data[88][135] = 0;
        pixel_data[88][136] = 0;
        pixel_data[88][137] = 0;
        pixel_data[88][138] = 0;
        pixel_data[88][139] = 0;
        pixel_data[88][140] = 0;
        pixel_data[88][141] = 0;
        pixel_data[88][142] = 0;
        pixel_data[88][143] = 0;
        pixel_data[88][144] = 0;
        pixel_data[88][145] = 0;
        pixel_data[88][146] = 0;
        pixel_data[88][147] = 0;
        pixel_data[88][148] = 0;
        pixel_data[88][149] = 0;
        pixel_data[88][150] = 0;
        pixel_data[88][151] = 0;
        pixel_data[88][152] = 0;
        pixel_data[88][153] = 0;
        pixel_data[88][154] = 0;
        pixel_data[88][155] = 0;
        pixel_data[88][156] = 0;
        pixel_data[88][157] = 0;
        pixel_data[88][158] = 0;
        pixel_data[88][159] = 0;
        pixel_data[88][160] = 0;
        pixel_data[88][161] = 0;
        pixel_data[88][162] = 0;
        pixel_data[88][163] = 0;
        pixel_data[88][164] = 0;
        pixel_data[88][165] = 0;
        pixel_data[88][166] = 0;
        pixel_data[88][167] = 0;
        pixel_data[88][168] = 0;
        pixel_data[88][169] = 0;
        pixel_data[88][170] = 0;
        pixel_data[88][171] = 0;
        pixel_data[88][172] = 0;
        pixel_data[88][173] = 0;
        pixel_data[88][174] = 0;
        pixel_data[88][175] = 0;
        pixel_data[88][176] = 0;
        pixel_data[88][177] = 0;
        pixel_data[88][178] = 0;
        pixel_data[88][179] = 0;
        pixel_data[88][180] = 0;
        pixel_data[88][181] = 0;
        pixel_data[88][182] = 0;
        pixel_data[88][183] = 0;
        pixel_data[88][184] = 0;
        pixel_data[88][185] = 0;
        pixel_data[88][186] = 0;
        pixel_data[88][187] = 0;
        pixel_data[88][188] = 0;
        pixel_data[88][189] = 0;
        pixel_data[88][190] = 0;
        pixel_data[88][191] = 0;
        pixel_data[88][192] = 0;
        pixel_data[88][193] = 0;
        pixel_data[88][194] = 0;
        pixel_data[88][195] = 0;
        pixel_data[88][196] = 0;
        pixel_data[88][197] = 0;
        pixel_data[88][198] = 0;
        pixel_data[88][199] = 0; // y=88
        pixel_data[89][0] = 0;
        pixel_data[89][1] = 0;
        pixel_data[89][2] = 0;
        pixel_data[89][3] = 0;
        pixel_data[89][4] = 0;
        pixel_data[89][5] = 0;
        pixel_data[89][6] = 0;
        pixel_data[89][7] = 0;
        pixel_data[89][8] = 0;
        pixel_data[89][9] = 0;
        pixel_data[89][10] = 0;
        pixel_data[89][11] = 0;
        pixel_data[89][12] = 0;
        pixel_data[89][13] = 0;
        pixel_data[89][14] = 0;
        pixel_data[89][15] = 0;
        pixel_data[89][16] = 0;
        pixel_data[89][17] = 0;
        pixel_data[89][18] = 0;
        pixel_data[89][19] = 0;
        pixel_data[89][20] = 0;
        pixel_data[89][21] = 0;
        pixel_data[89][22] = 0;
        pixel_data[89][23] = 0;
        pixel_data[89][24] = 0;
        pixel_data[89][25] = 0;
        pixel_data[89][26] = 0;
        pixel_data[89][27] = 0;
        pixel_data[89][28] = 0;
        pixel_data[89][29] = 0;
        pixel_data[89][30] = 0;
        pixel_data[89][31] = 0;
        pixel_data[89][32] = 0;
        pixel_data[89][33] = 0;
        pixel_data[89][34] = 0;
        pixel_data[89][35] = 0;
        pixel_data[89][36] = 0;
        pixel_data[89][37] = 0;
        pixel_data[89][38] = 0;
        pixel_data[89][39] = 0;
        pixel_data[89][40] = 0;
        pixel_data[89][41] = 0;
        pixel_data[89][42] = 0;
        pixel_data[89][43] = 0;
        pixel_data[89][44] = 0;
        pixel_data[89][45] = 0;
        pixel_data[89][46] = 0;
        pixel_data[89][47] = 0;
        pixel_data[89][48] = 0;
        pixel_data[89][49] = 0;
        pixel_data[89][50] = 0;
        pixel_data[89][51] = 0;
        pixel_data[89][52] = 0;
        pixel_data[89][53] = 0;
        pixel_data[89][54] = 0;
        pixel_data[89][55] = 0;
        pixel_data[89][56] = 0;
        pixel_data[89][57] = 0;
        pixel_data[89][58] = 0;
        pixel_data[89][59] = 0;
        pixel_data[89][60] = 0;
        pixel_data[89][61] = 0;
        pixel_data[89][62] = 0;
        pixel_data[89][63] = 0;
        pixel_data[89][64] = 0;
        pixel_data[89][65] = 0;
        pixel_data[89][66] = 0;
        pixel_data[89][67] = 0;
        pixel_data[89][68] = 0;
        pixel_data[89][69] = 0;
        pixel_data[89][70] = 0;
        pixel_data[89][71] = 0;
        pixel_data[89][72] = 0;
        pixel_data[89][73] = 0;
        pixel_data[89][74] = 0;
        pixel_data[89][75] = 0;
        pixel_data[89][76] = 0;
        pixel_data[89][77] = 0;
        pixel_data[89][78] = 0;
        pixel_data[89][79] = 0;
        pixel_data[89][80] = 0;
        pixel_data[89][81] = 0;
        pixel_data[89][82] = 0;
        pixel_data[89][83] = 0;
        pixel_data[89][84] = 0;
        pixel_data[89][85] = 0;
        pixel_data[89][86] = 0;
        pixel_data[89][87] = 0;
        pixel_data[89][88] = 0;
        pixel_data[89][89] = 0;
        pixel_data[89][90] = 0;
        pixel_data[89][91] = 0;
        pixel_data[89][92] = 0;
        pixel_data[89][93] = 0;
        pixel_data[89][94] = 0;
        pixel_data[89][95] = 0;
        pixel_data[89][96] = 0;
        pixel_data[89][97] = 0;
        pixel_data[89][98] = 0;
        pixel_data[89][99] = 0;
        pixel_data[89][100] = 0;
        pixel_data[89][101] = 0;
        pixel_data[89][102] = 0;
        pixel_data[89][103] = 0;
        pixel_data[89][104] = 0;
        pixel_data[89][105] = 0;
        pixel_data[89][106] = 0;
        pixel_data[89][107] = 0;
        pixel_data[89][108] = 0;
        pixel_data[89][109] = 0;
        pixel_data[89][110] = 0;
        pixel_data[89][111] = 0;
        pixel_data[89][112] = 0;
        pixel_data[89][113] = 0;
        pixel_data[89][114] = 0;
        pixel_data[89][115] = 0;
        pixel_data[89][116] = 0;
        pixel_data[89][117] = 0;
        pixel_data[89][118] = 0;
        pixel_data[89][119] = 0;
        pixel_data[89][120] = 0;
        pixel_data[89][121] = 0;
        pixel_data[89][122] = 0;
        pixel_data[89][123] = 0;
        pixel_data[89][124] = 0;
        pixel_data[89][125] = 0;
        pixel_data[89][126] = 0;
        pixel_data[89][127] = 0;
        pixel_data[89][128] = 0;
        pixel_data[89][129] = 0;
        pixel_data[89][130] = 0;
        pixel_data[89][131] = 0;
        pixel_data[89][132] = 0;
        pixel_data[89][133] = 0;
        pixel_data[89][134] = 0;
        pixel_data[89][135] = 0;
        pixel_data[89][136] = 0;
        pixel_data[89][137] = 0;
        pixel_data[89][138] = 0;
        pixel_data[89][139] = 0;
        pixel_data[89][140] = 0;
        pixel_data[89][141] = 0;
        pixel_data[89][142] = 0;
        pixel_data[89][143] = 0;
        pixel_data[89][144] = 0;
        pixel_data[89][145] = 0;
        pixel_data[89][146] = 0;
        pixel_data[89][147] = 0;
        pixel_data[89][148] = 0;
        pixel_data[89][149] = 0;
        pixel_data[89][150] = 0;
        pixel_data[89][151] = 0;
        pixel_data[89][152] = 0;
        pixel_data[89][153] = 0;
        pixel_data[89][154] = 0;
        pixel_data[89][155] = 0;
        pixel_data[89][156] = 0;
        pixel_data[89][157] = 0;
        pixel_data[89][158] = 0;
        pixel_data[89][159] = 0;
        pixel_data[89][160] = 0;
        pixel_data[89][161] = 0;
        pixel_data[89][162] = 0;
        pixel_data[89][163] = 0;
        pixel_data[89][164] = 0;
        pixel_data[89][165] = 0;
        pixel_data[89][166] = 0;
        pixel_data[89][167] = 0;
        pixel_data[89][168] = 0;
        pixel_data[89][169] = 0;
        pixel_data[89][170] = 0;
        pixel_data[89][171] = 0;
        pixel_data[89][172] = 0;
        pixel_data[89][173] = 0;
        pixel_data[89][174] = 0;
        pixel_data[89][175] = 0;
        pixel_data[89][176] = 0;
        pixel_data[89][177] = 0;
        pixel_data[89][178] = 0;
        pixel_data[89][179] = 0;
        pixel_data[89][180] = 0;
        pixel_data[89][181] = 0;
        pixel_data[89][182] = 0;
        pixel_data[89][183] = 0;
        pixel_data[89][184] = 0;
        pixel_data[89][185] = 0;
        pixel_data[89][186] = 0;
        pixel_data[89][187] = 0;
        pixel_data[89][188] = 0;
        pixel_data[89][189] = 0;
        pixel_data[89][190] = 0;
        pixel_data[89][191] = 0;
        pixel_data[89][192] = 0;
        pixel_data[89][193] = 0;
        pixel_data[89][194] = 0;
        pixel_data[89][195] = 0;
        pixel_data[89][196] = 0;
        pixel_data[89][197] = 0;
        pixel_data[89][198] = 0;
        pixel_data[89][199] = 0; // y=89
        pixel_data[90][0] = 0;
        pixel_data[90][1] = 0;
        pixel_data[90][2] = 0;
        pixel_data[90][3] = 0;
        pixel_data[90][4] = 0;
        pixel_data[90][5] = 0;
        pixel_data[90][6] = 0;
        pixel_data[90][7] = 0;
        pixel_data[90][8] = 0;
        pixel_data[90][9] = 0;
        pixel_data[90][10] = 0;
        pixel_data[90][11] = 0;
        pixel_data[90][12] = 0;
        pixel_data[90][13] = 0;
        pixel_data[90][14] = 0;
        pixel_data[90][15] = 0;
        pixel_data[90][16] = 0;
        pixel_data[90][17] = 0;
        pixel_data[90][18] = 0;
        pixel_data[90][19] = 0;
        pixel_data[90][20] = 0;
        pixel_data[90][21] = 0;
        pixel_data[90][22] = 0;
        pixel_data[90][23] = 0;
        pixel_data[90][24] = 0;
        pixel_data[90][25] = 0;
        pixel_data[90][26] = 0;
        pixel_data[90][27] = 0;
        pixel_data[90][28] = 0;
        pixel_data[90][29] = 0;
        pixel_data[90][30] = 0;
        pixel_data[90][31] = 0;
        pixel_data[90][32] = 0;
        pixel_data[90][33] = 0;
        pixel_data[90][34] = 0;
        pixel_data[90][35] = 0;
        pixel_data[90][36] = 0;
        pixel_data[90][37] = 0;
        pixel_data[90][38] = 0;
        pixel_data[90][39] = 0;
        pixel_data[90][40] = 0;
        pixel_data[90][41] = 0;
        pixel_data[90][42] = 0;
        pixel_data[90][43] = 0;
        pixel_data[90][44] = 0;
        pixel_data[90][45] = 0;
        pixel_data[90][46] = 0;
        pixel_data[90][47] = 0;
        pixel_data[90][48] = 0;
        pixel_data[90][49] = 0;
        pixel_data[90][50] = 0;
        pixel_data[90][51] = 0;
        pixel_data[90][52] = 0;
        pixel_data[90][53] = 0;
        pixel_data[90][54] = 0;
        pixel_data[90][55] = 0;
        pixel_data[90][56] = 0;
        pixel_data[90][57] = 0;
        pixel_data[90][58] = 0;
        pixel_data[90][59] = 0;
        pixel_data[90][60] = 0;
        pixel_data[90][61] = 0;
        pixel_data[90][62] = 0;
        pixel_data[90][63] = 0;
        pixel_data[90][64] = 0;
        pixel_data[90][65] = 0;
        pixel_data[90][66] = 0;
        pixel_data[90][67] = 0;
        pixel_data[90][68] = 0;
        pixel_data[90][69] = 0;
        pixel_data[90][70] = 0;
        pixel_data[90][71] = 0;
        pixel_data[90][72] = 0;
        pixel_data[90][73] = 0;
        pixel_data[90][74] = 0;
        pixel_data[90][75] = 0;
        pixel_data[90][76] = 0;
        pixel_data[90][77] = 0;
        pixel_data[90][78] = 0;
        pixel_data[90][79] = 0;
        pixel_data[90][80] = 0;
        pixel_data[90][81] = 0;
        pixel_data[90][82] = 0;
        pixel_data[90][83] = 0;
        pixel_data[90][84] = 0;
        pixel_data[90][85] = 0;
        pixel_data[90][86] = 0;
        pixel_data[90][87] = 0;
        pixel_data[90][88] = 0;
        pixel_data[90][89] = 0;
        pixel_data[90][90] = 0;
        pixel_data[90][91] = 0;
        pixel_data[90][92] = 0;
        pixel_data[90][93] = 0;
        pixel_data[90][94] = 0;
        pixel_data[90][95] = 0;
        pixel_data[90][96] = 0;
        pixel_data[90][97] = 0;
        pixel_data[90][98] = 0;
        pixel_data[90][99] = 0;
        pixel_data[90][100] = 0;
        pixel_data[90][101] = 0;
        pixel_data[90][102] = 0;
        pixel_data[90][103] = 0;
        pixel_data[90][104] = 0;
        pixel_data[90][105] = 0;
        pixel_data[90][106] = 0;
        pixel_data[90][107] = 0;
        pixel_data[90][108] = 0;
        pixel_data[90][109] = 0;
        pixel_data[90][110] = 0;
        pixel_data[90][111] = 0;
        pixel_data[90][112] = 0;
        pixel_data[90][113] = 0;
        pixel_data[90][114] = 0;
        pixel_data[90][115] = 0;
        pixel_data[90][116] = 0;
        pixel_data[90][117] = 0;
        pixel_data[90][118] = 0;
        pixel_data[90][119] = 0;
        pixel_data[90][120] = 0;
        pixel_data[90][121] = 0;
        pixel_data[90][122] = 0;
        pixel_data[90][123] = 0;
        pixel_data[90][124] = 0;
        pixel_data[90][125] = 0;
        pixel_data[90][126] = 0;
        pixel_data[90][127] = 0;
        pixel_data[90][128] = 0;
        pixel_data[90][129] = 0;
        pixel_data[90][130] = 0;
        pixel_data[90][131] = 0;
        pixel_data[90][132] = 0;
        pixel_data[90][133] = 0;
        pixel_data[90][134] = 0;
        pixel_data[90][135] = 0;
        pixel_data[90][136] = 0;
        pixel_data[90][137] = 0;
        pixel_data[90][138] = 0;
        pixel_data[90][139] = 0;
        pixel_data[90][140] = 0;
        pixel_data[90][141] = 0;
        pixel_data[90][142] = 0;
        pixel_data[90][143] = 0;
        pixel_data[90][144] = 0;
        pixel_data[90][145] = 0;
        pixel_data[90][146] = 0;
        pixel_data[90][147] = 0;
        pixel_data[90][148] = 0;
        pixel_data[90][149] = 0;
        pixel_data[90][150] = 0;
        pixel_data[90][151] = 0;
        pixel_data[90][152] = 0;
        pixel_data[90][153] = 0;
        pixel_data[90][154] = 0;
        pixel_data[90][155] = 0;
        pixel_data[90][156] = 0;
        pixel_data[90][157] = 0;
        pixel_data[90][158] = 0;
        pixel_data[90][159] = 0;
        pixel_data[90][160] = 0;
        pixel_data[90][161] = 0;
        pixel_data[90][162] = 0;
        pixel_data[90][163] = 0;
        pixel_data[90][164] = 0;
        pixel_data[90][165] = 0;
        pixel_data[90][166] = 0;
        pixel_data[90][167] = 0;
        pixel_data[90][168] = 0;
        pixel_data[90][169] = 0;
        pixel_data[90][170] = 0;
        pixel_data[90][171] = 0;
        pixel_data[90][172] = 0;
        pixel_data[90][173] = 0;
        pixel_data[90][174] = 0;
        pixel_data[90][175] = 0;
        pixel_data[90][176] = 0;
        pixel_data[90][177] = 0;
        pixel_data[90][178] = 0;
        pixel_data[90][179] = 0;
        pixel_data[90][180] = 0;
        pixel_data[90][181] = 0;
        pixel_data[90][182] = 0;
        pixel_data[90][183] = 0;
        pixel_data[90][184] = 0;
        pixel_data[90][185] = 0;
        pixel_data[90][186] = 0;
        pixel_data[90][187] = 0;
        pixel_data[90][188] = 0;
        pixel_data[90][189] = 0;
        pixel_data[90][190] = 0;
        pixel_data[90][191] = 0;
        pixel_data[90][192] = 0;
        pixel_data[90][193] = 0;
        pixel_data[90][194] = 0;
        pixel_data[90][195] = 0;
        pixel_data[90][196] = 0;
        pixel_data[90][197] = 0;
        pixel_data[90][198] = 0;
        pixel_data[90][199] = 0; // y=90
        pixel_data[91][0] = 0;
        pixel_data[91][1] = 0;
        pixel_data[91][2] = 0;
        pixel_data[91][3] = 0;
        pixel_data[91][4] = 0;
        pixel_data[91][5] = 0;
        pixel_data[91][6] = 0;
        pixel_data[91][7] = 0;
        pixel_data[91][8] = 0;
        pixel_data[91][9] = 0;
        pixel_data[91][10] = 0;
        pixel_data[91][11] = 0;
        pixel_data[91][12] = 0;
        pixel_data[91][13] = 0;
        pixel_data[91][14] = 0;
        pixel_data[91][15] = 0;
        pixel_data[91][16] = 0;
        pixel_data[91][17] = 0;
        pixel_data[91][18] = 0;
        pixel_data[91][19] = 0;
        pixel_data[91][20] = 0;
        pixel_data[91][21] = 0;
        pixel_data[91][22] = 0;
        pixel_data[91][23] = 0;
        pixel_data[91][24] = 0;
        pixel_data[91][25] = 0;
        pixel_data[91][26] = 0;
        pixel_data[91][27] = 0;
        pixel_data[91][28] = 0;
        pixel_data[91][29] = 0;
        pixel_data[91][30] = 0;
        pixel_data[91][31] = 0;
        pixel_data[91][32] = 0;
        pixel_data[91][33] = 0;
        pixel_data[91][34] = 0;
        pixel_data[91][35] = 0;
        pixel_data[91][36] = 0;
        pixel_data[91][37] = 0;
        pixel_data[91][38] = 0;
        pixel_data[91][39] = 0;
        pixel_data[91][40] = 0;
        pixel_data[91][41] = 0;
        pixel_data[91][42] = 0;
        pixel_data[91][43] = 0;
        pixel_data[91][44] = 0;
        pixel_data[91][45] = 0;
        pixel_data[91][46] = 0;
        pixel_data[91][47] = 0;
        pixel_data[91][48] = 0;
        pixel_data[91][49] = 0;
        pixel_data[91][50] = 0;
        pixel_data[91][51] = 0;
        pixel_data[91][52] = 0;
        pixel_data[91][53] = 0;
        pixel_data[91][54] = 0;
        pixel_data[91][55] = 0;
        pixel_data[91][56] = 0;
        pixel_data[91][57] = 0;
        pixel_data[91][58] = 0;
        pixel_data[91][59] = 0;
        pixel_data[91][60] = 0;
        pixel_data[91][61] = 0;
        pixel_data[91][62] = 0;
        pixel_data[91][63] = 0;
        pixel_data[91][64] = 0;
        pixel_data[91][65] = 0;
        pixel_data[91][66] = 0;
        pixel_data[91][67] = 0;
        pixel_data[91][68] = 0;
        pixel_data[91][69] = 0;
        pixel_data[91][70] = 0;
        pixel_data[91][71] = 0;
        pixel_data[91][72] = 0;
        pixel_data[91][73] = 0;
        pixel_data[91][74] = 0;
        pixel_data[91][75] = 0;
        pixel_data[91][76] = 0;
        pixel_data[91][77] = 0;
        pixel_data[91][78] = 0;
        pixel_data[91][79] = 0;
        pixel_data[91][80] = 0;
        pixel_data[91][81] = 0;
        pixel_data[91][82] = 0;
        pixel_data[91][83] = 0;
        pixel_data[91][84] = 0;
        pixel_data[91][85] = 0;
        pixel_data[91][86] = 0;
        pixel_data[91][87] = 0;
        pixel_data[91][88] = 0;
        pixel_data[91][89] = 0;
        pixel_data[91][90] = 0;
        pixel_data[91][91] = 0;
        pixel_data[91][92] = 0;
        pixel_data[91][93] = 0;
        pixel_data[91][94] = 0;
        pixel_data[91][95] = 0;
        pixel_data[91][96] = 0;
        pixel_data[91][97] = 0;
        pixel_data[91][98] = 0;
        pixel_data[91][99] = 0;
        pixel_data[91][100] = 0;
        pixel_data[91][101] = 0;
        pixel_data[91][102] = 0;
        pixel_data[91][103] = 0;
        pixel_data[91][104] = 0;
        pixel_data[91][105] = 0;
        pixel_data[91][106] = 0;
        pixel_data[91][107] = 0;
        pixel_data[91][108] = 0;
        pixel_data[91][109] = 0;
        pixel_data[91][110] = 0;
        pixel_data[91][111] = 0;
        pixel_data[91][112] = 0;
        pixel_data[91][113] = 0;
        pixel_data[91][114] = 0;
        pixel_data[91][115] = 0;
        pixel_data[91][116] = 0;
        pixel_data[91][117] = 0;
        pixel_data[91][118] = 0;
        pixel_data[91][119] = 0;
        pixel_data[91][120] = 0;
        pixel_data[91][121] = 0;
        pixel_data[91][122] = 0;
        pixel_data[91][123] = 0;
        pixel_data[91][124] = 0;
        pixel_data[91][125] = 0;
        pixel_data[91][126] = 0;
        pixel_data[91][127] = 0;
        pixel_data[91][128] = 0;
        pixel_data[91][129] = 0;
        pixel_data[91][130] = 0;
        pixel_data[91][131] = 0;
        pixel_data[91][132] = 0;
        pixel_data[91][133] = 0;
        pixel_data[91][134] = 0;
        pixel_data[91][135] = 0;
        pixel_data[91][136] = 0;
        pixel_data[91][137] = 0;
        pixel_data[91][138] = 0;
        pixel_data[91][139] = 0;
        pixel_data[91][140] = 0;
        pixel_data[91][141] = 0;
        pixel_data[91][142] = 0;
        pixel_data[91][143] = 0;
        pixel_data[91][144] = 0;
        pixel_data[91][145] = 0;
        pixel_data[91][146] = 0;
        pixel_data[91][147] = 0;
        pixel_data[91][148] = 0;
        pixel_data[91][149] = 0;
        pixel_data[91][150] = 0;
        pixel_data[91][151] = 0;
        pixel_data[91][152] = 0;
        pixel_data[91][153] = 0;
        pixel_data[91][154] = 0;
        pixel_data[91][155] = 0;
        pixel_data[91][156] = 0;
        pixel_data[91][157] = 0;
        pixel_data[91][158] = 0;
        pixel_data[91][159] = 0;
        pixel_data[91][160] = 0;
        pixel_data[91][161] = 0;
        pixel_data[91][162] = 0;
        pixel_data[91][163] = 0;
        pixel_data[91][164] = 0;
        pixel_data[91][165] = 0;
        pixel_data[91][166] = 0;
        pixel_data[91][167] = 0;
        pixel_data[91][168] = 0;
        pixel_data[91][169] = 0;
        pixel_data[91][170] = 0;
        pixel_data[91][171] = 0;
        pixel_data[91][172] = 0;
        pixel_data[91][173] = 0;
        pixel_data[91][174] = 0;
        pixel_data[91][175] = 0;
        pixel_data[91][176] = 0;
        pixel_data[91][177] = 0;
        pixel_data[91][178] = 0;
        pixel_data[91][179] = 0;
        pixel_data[91][180] = 0;
        pixel_data[91][181] = 0;
        pixel_data[91][182] = 0;
        pixel_data[91][183] = 0;
        pixel_data[91][184] = 0;
        pixel_data[91][185] = 0;
        pixel_data[91][186] = 0;
        pixel_data[91][187] = 0;
        pixel_data[91][188] = 0;
        pixel_data[91][189] = 0;
        pixel_data[91][190] = 0;
        pixel_data[91][191] = 0;
        pixel_data[91][192] = 0;
        pixel_data[91][193] = 0;
        pixel_data[91][194] = 0;
        pixel_data[91][195] = 0;
        pixel_data[91][196] = 0;
        pixel_data[91][197] = 0;
        pixel_data[91][198] = 0;
        pixel_data[91][199] = 0; // y=91
        pixel_data[92][0] = 0;
        pixel_data[92][1] = 0;
        pixel_data[92][2] = 0;
        pixel_data[92][3] = 0;
        pixel_data[92][4] = 0;
        pixel_data[92][5] = 0;
        pixel_data[92][6] = 0;
        pixel_data[92][7] = 0;
        pixel_data[92][8] = 0;
        pixel_data[92][9] = 0;
        pixel_data[92][10] = 0;
        pixel_data[92][11] = 0;
        pixel_data[92][12] = 0;
        pixel_data[92][13] = 0;
        pixel_data[92][14] = 0;
        pixel_data[92][15] = 0;
        pixel_data[92][16] = 0;
        pixel_data[92][17] = 0;
        pixel_data[92][18] = 0;
        pixel_data[92][19] = 0;
        pixel_data[92][20] = 0;
        pixel_data[92][21] = 0;
        pixel_data[92][22] = 0;
        pixel_data[92][23] = 0;
        pixel_data[92][24] = 0;
        pixel_data[92][25] = 0;
        pixel_data[92][26] = 0;
        pixel_data[92][27] = 0;
        pixel_data[92][28] = 0;
        pixel_data[92][29] = 0;
        pixel_data[92][30] = 0;
        pixel_data[92][31] = 0;
        pixel_data[92][32] = 0;
        pixel_data[92][33] = 0;
        pixel_data[92][34] = 0;
        pixel_data[92][35] = 0;
        pixel_data[92][36] = 0;
        pixel_data[92][37] = 0;
        pixel_data[92][38] = 0;
        pixel_data[92][39] = 0;
        pixel_data[92][40] = 0;
        pixel_data[92][41] = 0;
        pixel_data[92][42] = 0;
        pixel_data[92][43] = 0;
        pixel_data[92][44] = 0;
        pixel_data[92][45] = 0;
        pixel_data[92][46] = 0;
        pixel_data[92][47] = 0;
        pixel_data[92][48] = 0;
        pixel_data[92][49] = 0;
        pixel_data[92][50] = 0;
        pixel_data[92][51] = 0;
        pixel_data[92][52] = 0;
        pixel_data[92][53] = 0;
        pixel_data[92][54] = 0;
        pixel_data[92][55] = 0;
        pixel_data[92][56] = 0;
        pixel_data[92][57] = 0;
        pixel_data[92][58] = 0;
        pixel_data[92][59] = 0;
        pixel_data[92][60] = 0;
        pixel_data[92][61] = 0;
        pixel_data[92][62] = 0;
        pixel_data[92][63] = 0;
        pixel_data[92][64] = 0;
        pixel_data[92][65] = 0;
        pixel_data[92][66] = 0;
        pixel_data[92][67] = 0;
        pixel_data[92][68] = 0;
        pixel_data[92][69] = 0;
        pixel_data[92][70] = 0;
        pixel_data[92][71] = 0;
        pixel_data[92][72] = 0;
        pixel_data[92][73] = 0;
        pixel_data[92][74] = 0;
        pixel_data[92][75] = 0;
        pixel_data[92][76] = 0;
        pixel_data[92][77] = 0;
        pixel_data[92][78] = 0;
        pixel_data[92][79] = 0;
        pixel_data[92][80] = 0;
        pixel_data[92][81] = 0;
        pixel_data[92][82] = 0;
        pixel_data[92][83] = 0;
        pixel_data[92][84] = 0;
        pixel_data[92][85] = 0;
        pixel_data[92][86] = 0;
        pixel_data[92][87] = 0;
        pixel_data[92][88] = 0;
        pixel_data[92][89] = 0;
        pixel_data[92][90] = 0;
        pixel_data[92][91] = 0;
        pixel_data[92][92] = 0;
        pixel_data[92][93] = 0;
        pixel_data[92][94] = 0;
        pixel_data[92][95] = 0;
        pixel_data[92][96] = 0;
        pixel_data[92][97] = 0;
        pixel_data[92][98] = 0;
        pixel_data[92][99] = 0;
        pixel_data[92][100] = 0;
        pixel_data[92][101] = 0;
        pixel_data[92][102] = 0;
        pixel_data[92][103] = 0;
        pixel_data[92][104] = 0;
        pixel_data[92][105] = 0;
        pixel_data[92][106] = 0;
        pixel_data[92][107] = 0;
        pixel_data[92][108] = 0;
        pixel_data[92][109] = 0;
        pixel_data[92][110] = 0;
        pixel_data[92][111] = 0;
        pixel_data[92][112] = 0;
        pixel_data[92][113] = 0;
        pixel_data[92][114] = 0;
        pixel_data[92][115] = 0;
        pixel_data[92][116] = 0;
        pixel_data[92][117] = 0;
        pixel_data[92][118] = 0;
        pixel_data[92][119] = 0;
        pixel_data[92][120] = 0;
        pixel_data[92][121] = 0;
        pixel_data[92][122] = 0;
        pixel_data[92][123] = 0;
        pixel_data[92][124] = 0;
        pixel_data[92][125] = 0;
        pixel_data[92][126] = 0;
        pixel_data[92][127] = 0;
        pixel_data[92][128] = 0;
        pixel_data[92][129] = 0;
        pixel_data[92][130] = 0;
        pixel_data[92][131] = 0;
        pixel_data[92][132] = 0;
        pixel_data[92][133] = 0;
        pixel_data[92][134] = 0;
        pixel_data[92][135] = 0;
        pixel_data[92][136] = 0;
        pixel_data[92][137] = 0;
        pixel_data[92][138] = 0;
        pixel_data[92][139] = 0;
        pixel_data[92][140] = 0;
        pixel_data[92][141] = 0;
        pixel_data[92][142] = 0;
        pixel_data[92][143] = 0;
        pixel_data[92][144] = 0;
        pixel_data[92][145] = 0;
        pixel_data[92][146] = 0;
        pixel_data[92][147] = 0;
        pixel_data[92][148] = 0;
        pixel_data[92][149] = 0;
        pixel_data[92][150] = 0;
        pixel_data[92][151] = 0;
        pixel_data[92][152] = 0;
        pixel_data[92][153] = 0;
        pixel_data[92][154] = 0;
        pixel_data[92][155] = 0;
        pixel_data[92][156] = 0;
        pixel_data[92][157] = 0;
        pixel_data[92][158] = 0;
        pixel_data[92][159] = 0;
        pixel_data[92][160] = 0;
        pixel_data[92][161] = 0;
        pixel_data[92][162] = 0;
        pixel_data[92][163] = 0;
        pixel_data[92][164] = 0;
        pixel_data[92][165] = 0;
        pixel_data[92][166] = 0;
        pixel_data[92][167] = 0;
        pixel_data[92][168] = 0;
        pixel_data[92][169] = 0;
        pixel_data[92][170] = 0;
        pixel_data[92][171] = 0;
        pixel_data[92][172] = 0;
        pixel_data[92][173] = 0;
        pixel_data[92][174] = 0;
        pixel_data[92][175] = 0;
        pixel_data[92][176] = 0;
        pixel_data[92][177] = 0;
        pixel_data[92][178] = 0;
        pixel_data[92][179] = 0;
        pixel_data[92][180] = 0;
        pixel_data[92][181] = 0;
        pixel_data[92][182] = 0;
        pixel_data[92][183] = 0;
        pixel_data[92][184] = 0;
        pixel_data[92][185] = 0;
        pixel_data[92][186] = 0;
        pixel_data[92][187] = 0;
        pixel_data[92][188] = 0;
        pixel_data[92][189] = 0;
        pixel_data[92][190] = 0;
        pixel_data[92][191] = 0;
        pixel_data[92][192] = 0;
        pixel_data[92][193] = 0;
        pixel_data[92][194] = 0;
        pixel_data[92][195] = 0;
        pixel_data[92][196] = 0;
        pixel_data[92][197] = 0;
        pixel_data[92][198] = 0;
        pixel_data[92][199] = 0; // y=92
        pixel_data[93][0] = 0;
        pixel_data[93][1] = 0;
        pixel_data[93][2] = 0;
        pixel_data[93][3] = 0;
        pixel_data[93][4] = 0;
        pixel_data[93][5] = 0;
        pixel_data[93][6] = 0;
        pixel_data[93][7] = 0;
        pixel_data[93][8] = 0;
        pixel_data[93][9] = 0;
        pixel_data[93][10] = 0;
        pixel_data[93][11] = 0;
        pixel_data[93][12] = 0;
        pixel_data[93][13] = 0;
        pixel_data[93][14] = 0;
        pixel_data[93][15] = 0;
        pixel_data[93][16] = 0;
        pixel_data[93][17] = 0;
        pixel_data[93][18] = 0;
        pixel_data[93][19] = 0;
        pixel_data[93][20] = 0;
        pixel_data[93][21] = 0;
        pixel_data[93][22] = 0;
        pixel_data[93][23] = 0;
        pixel_data[93][24] = 0;
        pixel_data[93][25] = 0;
        pixel_data[93][26] = 0;
        pixel_data[93][27] = 0;
        pixel_data[93][28] = 0;
        pixel_data[93][29] = 0;
        pixel_data[93][30] = 0;
        pixel_data[93][31] = 0;
        pixel_data[93][32] = 0;
        pixel_data[93][33] = 0;
        pixel_data[93][34] = 0;
        pixel_data[93][35] = 0;
        pixel_data[93][36] = 0;
        pixel_data[93][37] = 0;
        pixel_data[93][38] = 0;
        pixel_data[93][39] = 0;
        pixel_data[93][40] = 0;
        pixel_data[93][41] = 0;
        pixel_data[93][42] = 0;
        pixel_data[93][43] = 0;
        pixel_data[93][44] = 0;
        pixel_data[93][45] = 0;
        pixel_data[93][46] = 0;
        pixel_data[93][47] = 0;
        pixel_data[93][48] = 0;
        pixel_data[93][49] = 0;
        pixel_data[93][50] = 0;
        pixel_data[93][51] = 0;
        pixel_data[93][52] = 0;
        pixel_data[93][53] = 0;
        pixel_data[93][54] = 0;
        pixel_data[93][55] = 0;
        pixel_data[93][56] = 0;
        pixel_data[93][57] = 0;
        pixel_data[93][58] = 0;
        pixel_data[93][59] = 0;
        pixel_data[93][60] = 0;
        pixel_data[93][61] = 0;
        pixel_data[93][62] = 0;
        pixel_data[93][63] = 0;
        pixel_data[93][64] = 0;
        pixel_data[93][65] = 0;
        pixel_data[93][66] = 0;
        pixel_data[93][67] = 0;
        pixel_data[93][68] = 0;
        pixel_data[93][69] = 0;
        pixel_data[93][70] = 0;
        pixel_data[93][71] = 0;
        pixel_data[93][72] = 0;
        pixel_data[93][73] = 0;
        pixel_data[93][74] = 0;
        pixel_data[93][75] = 0;
        pixel_data[93][76] = 0;
        pixel_data[93][77] = 0;
        pixel_data[93][78] = 0;
        pixel_data[93][79] = 0;
        pixel_data[93][80] = 0;
        pixel_data[93][81] = 0;
        pixel_data[93][82] = 0;
        pixel_data[93][83] = 0;
        pixel_data[93][84] = 0;
        pixel_data[93][85] = 0;
        pixel_data[93][86] = 0;
        pixel_data[93][87] = 0;
        pixel_data[93][88] = 0;
        pixel_data[93][89] = 0;
        pixel_data[93][90] = 0;
        pixel_data[93][91] = 0;
        pixel_data[93][92] = 0;
        pixel_data[93][93] = 0;
        pixel_data[93][94] = 0;
        pixel_data[93][95] = 0;
        pixel_data[93][96] = 0;
        pixel_data[93][97] = 0;
        pixel_data[93][98] = 0;
        pixel_data[93][99] = 0;
        pixel_data[93][100] = 0;
        pixel_data[93][101] = 0;
        pixel_data[93][102] = 0;
        pixel_data[93][103] = 0;
        pixel_data[93][104] = 0;
        pixel_data[93][105] = 0;
        pixel_data[93][106] = 0;
        pixel_data[93][107] = 0;
        pixel_data[93][108] = 0;
        pixel_data[93][109] = 0;
        pixel_data[93][110] = 0;
        pixel_data[93][111] = 0;
        pixel_data[93][112] = 0;
        pixel_data[93][113] = 0;
        pixel_data[93][114] = 0;
        pixel_data[93][115] = 0;
        pixel_data[93][116] = 0;
        pixel_data[93][117] = 0;
        pixel_data[93][118] = 0;
        pixel_data[93][119] = 0;
        pixel_data[93][120] = 0;
        pixel_data[93][121] = 0;
        pixel_data[93][122] = 0;
        pixel_data[93][123] = 0;
        pixel_data[93][124] = 0;
        pixel_data[93][125] = 0;
        pixel_data[93][126] = 0;
        pixel_data[93][127] = 0;
        pixel_data[93][128] = 0;
        pixel_data[93][129] = 0;
        pixel_data[93][130] = 0;
        pixel_data[93][131] = 0;
        pixel_data[93][132] = 0;
        pixel_data[93][133] = 0;
        pixel_data[93][134] = 0;
        pixel_data[93][135] = 0;
        pixel_data[93][136] = 0;
        pixel_data[93][137] = 0;
        pixel_data[93][138] = 0;
        pixel_data[93][139] = 0;
        pixel_data[93][140] = 0;
        pixel_data[93][141] = 0;
        pixel_data[93][142] = 0;
        pixel_data[93][143] = 0;
        pixel_data[93][144] = 0;
        pixel_data[93][145] = 0;
        pixel_data[93][146] = 0;
        pixel_data[93][147] = 0;
        pixel_data[93][148] = 0;
        pixel_data[93][149] = 0;
        pixel_data[93][150] = 0;
        pixel_data[93][151] = 0;
        pixel_data[93][152] = 0;
        pixel_data[93][153] = 0;
        pixel_data[93][154] = 0;
        pixel_data[93][155] = 0;
        pixel_data[93][156] = 0;
        pixel_data[93][157] = 0;
        pixel_data[93][158] = 0;
        pixel_data[93][159] = 0;
        pixel_data[93][160] = 0;
        pixel_data[93][161] = 0;
        pixel_data[93][162] = 0;
        pixel_data[93][163] = 0;
        pixel_data[93][164] = 0;
        pixel_data[93][165] = 0;
        pixel_data[93][166] = 0;
        pixel_data[93][167] = 0;
        pixel_data[93][168] = 0;
        pixel_data[93][169] = 0;
        pixel_data[93][170] = 0;
        pixel_data[93][171] = 0;
        pixel_data[93][172] = 0;
        pixel_data[93][173] = 0;
        pixel_data[93][174] = 0;
        pixel_data[93][175] = 0;
        pixel_data[93][176] = 0;
        pixel_data[93][177] = 0;
        pixel_data[93][178] = 0;
        pixel_data[93][179] = 0;
        pixel_data[93][180] = 0;
        pixel_data[93][181] = 0;
        pixel_data[93][182] = 0;
        pixel_data[93][183] = 0;
        pixel_data[93][184] = 0;
        pixel_data[93][185] = 0;
        pixel_data[93][186] = 0;
        pixel_data[93][187] = 0;
        pixel_data[93][188] = 0;
        pixel_data[93][189] = 0;
        pixel_data[93][190] = 0;
        pixel_data[93][191] = 0;
        pixel_data[93][192] = 0;
        pixel_data[93][193] = 0;
        pixel_data[93][194] = 0;
        pixel_data[93][195] = 0;
        pixel_data[93][196] = 0;
        pixel_data[93][197] = 0;
        pixel_data[93][198] = 0;
        pixel_data[93][199] = 0; // y=93
        pixel_data[94][0] = 0;
        pixel_data[94][1] = 0;
        pixel_data[94][2] = 0;
        pixel_data[94][3] = 0;
        pixel_data[94][4] = 0;
        pixel_data[94][5] = 0;
        pixel_data[94][6] = 0;
        pixel_data[94][7] = 0;
        pixel_data[94][8] = 0;
        pixel_data[94][9] = 0;
        pixel_data[94][10] = 0;
        pixel_data[94][11] = 0;
        pixel_data[94][12] = 0;
        pixel_data[94][13] = 0;
        pixel_data[94][14] = 0;
        pixel_data[94][15] = 0;
        pixel_data[94][16] = 0;
        pixel_data[94][17] = 0;
        pixel_data[94][18] = 0;
        pixel_data[94][19] = 0;
        pixel_data[94][20] = 0;
        pixel_data[94][21] = 0;
        pixel_data[94][22] = 0;
        pixel_data[94][23] = 0;
        pixel_data[94][24] = 0;
        pixel_data[94][25] = 0;
        pixel_data[94][26] = 0;
        pixel_data[94][27] = 0;
        pixel_data[94][28] = 0;
        pixel_data[94][29] = 0;
        pixel_data[94][30] = 0;
        pixel_data[94][31] = 0;
        pixel_data[94][32] = 0;
        pixel_data[94][33] = 0;
        pixel_data[94][34] = 0;
        pixel_data[94][35] = 0;
        pixel_data[94][36] = 0;
        pixel_data[94][37] = 0;
        pixel_data[94][38] = 0;
        pixel_data[94][39] = 0;
        pixel_data[94][40] = 0;
        pixel_data[94][41] = 0;
        pixel_data[94][42] = 0;
        pixel_data[94][43] = 0;
        pixel_data[94][44] = 0;
        pixel_data[94][45] = 0;
        pixel_data[94][46] = 0;
        pixel_data[94][47] = 0;
        pixel_data[94][48] = 0;
        pixel_data[94][49] = 0;
        pixel_data[94][50] = 0;
        pixel_data[94][51] = 0;
        pixel_data[94][52] = 0;
        pixel_data[94][53] = 0;
        pixel_data[94][54] = 0;
        pixel_data[94][55] = 0;
        pixel_data[94][56] = 0;
        pixel_data[94][57] = 0;
        pixel_data[94][58] = 0;
        pixel_data[94][59] = 0;
        pixel_data[94][60] = 0;
        pixel_data[94][61] = 0;
        pixel_data[94][62] = 0;
        pixel_data[94][63] = 0;
        pixel_data[94][64] = 0;
        pixel_data[94][65] = 0;
        pixel_data[94][66] = 0;
        pixel_data[94][67] = 0;
        pixel_data[94][68] = 0;
        pixel_data[94][69] = 0;
        pixel_data[94][70] = 0;
        pixel_data[94][71] = 0;
        pixel_data[94][72] = 0;
        pixel_data[94][73] = 0;
        pixel_data[94][74] = 0;
        pixel_data[94][75] = 0;
        pixel_data[94][76] = 0;
        pixel_data[94][77] = 0;
        pixel_data[94][78] = 0;
        pixel_data[94][79] = 0;
        pixel_data[94][80] = 0;
        pixel_data[94][81] = 0;
        pixel_data[94][82] = 0;
        pixel_data[94][83] = 0;
        pixel_data[94][84] = 0;
        pixel_data[94][85] = 0;
        pixel_data[94][86] = 0;
        pixel_data[94][87] = 0;
        pixel_data[94][88] = 0;
        pixel_data[94][89] = 0;
        pixel_data[94][90] = 0;
        pixel_data[94][91] = 0;
        pixel_data[94][92] = 0;
        pixel_data[94][93] = 0;
        pixel_data[94][94] = 0;
        pixel_data[94][95] = 0;
        pixel_data[94][96] = 0;
        pixel_data[94][97] = 0;
        pixel_data[94][98] = 0;
        pixel_data[94][99] = 0;
        pixel_data[94][100] = 0;
        pixel_data[94][101] = 0;
        pixel_data[94][102] = 0;
        pixel_data[94][103] = 0;
        pixel_data[94][104] = 0;
        pixel_data[94][105] = 0;
        pixel_data[94][106] = 0;
        pixel_data[94][107] = 0;
        pixel_data[94][108] = 0;
        pixel_data[94][109] = 0;
        pixel_data[94][110] = 0;
        pixel_data[94][111] = 0;
        pixel_data[94][112] = 0;
        pixel_data[94][113] = 0;
        pixel_data[94][114] = 0;
        pixel_data[94][115] = 0;
        pixel_data[94][116] = 0;
        pixel_data[94][117] = 0;
        pixel_data[94][118] = 0;
        pixel_data[94][119] = 0;
        pixel_data[94][120] = 0;
        pixel_data[94][121] = 0;
        pixel_data[94][122] = 0;
        pixel_data[94][123] = 0;
        pixel_data[94][124] = 0;
        pixel_data[94][125] = 0;
        pixel_data[94][126] = 0;
        pixel_data[94][127] = 0;
        pixel_data[94][128] = 0;
        pixel_data[94][129] = 0;
        pixel_data[94][130] = 0;
        pixel_data[94][131] = 0;
        pixel_data[94][132] = 0;
        pixel_data[94][133] = 0;
        pixel_data[94][134] = 0;
        pixel_data[94][135] = 0;
        pixel_data[94][136] = 0;
        pixel_data[94][137] = 0;
        pixel_data[94][138] = 0;
        pixel_data[94][139] = 0;
        pixel_data[94][140] = 0;
        pixel_data[94][141] = 0;
        pixel_data[94][142] = 0;
        pixel_data[94][143] = 0;
        pixel_data[94][144] = 0;
        pixel_data[94][145] = 0;
        pixel_data[94][146] = 0;
        pixel_data[94][147] = 0;
        pixel_data[94][148] = 0;
        pixel_data[94][149] = 0;
        pixel_data[94][150] = 0;
        pixel_data[94][151] = 0;
        pixel_data[94][152] = 0;
        pixel_data[94][153] = 0;
        pixel_data[94][154] = 0;
        pixel_data[94][155] = 0;
        pixel_data[94][156] = 0;
        pixel_data[94][157] = 0;
        pixel_data[94][158] = 0;
        pixel_data[94][159] = 0;
        pixel_data[94][160] = 0;
        pixel_data[94][161] = 0;
        pixel_data[94][162] = 0;
        pixel_data[94][163] = 0;
        pixel_data[94][164] = 0;
        pixel_data[94][165] = 0;
        pixel_data[94][166] = 0;
        pixel_data[94][167] = 0;
        pixel_data[94][168] = 0;
        pixel_data[94][169] = 0;
        pixel_data[94][170] = 0;
        pixel_data[94][171] = 0;
        pixel_data[94][172] = 0;
        pixel_data[94][173] = 0;
        pixel_data[94][174] = 0;
        pixel_data[94][175] = 0;
        pixel_data[94][176] = 0;
        pixel_data[94][177] = 0;
        pixel_data[94][178] = 0;
        pixel_data[94][179] = 0;
        pixel_data[94][180] = 0;
        pixel_data[94][181] = 0;
        pixel_data[94][182] = 0;
        pixel_data[94][183] = 0;
        pixel_data[94][184] = 0;
        pixel_data[94][185] = 0;
        pixel_data[94][186] = 0;
        pixel_data[94][187] = 0;
        pixel_data[94][188] = 0;
        pixel_data[94][189] = 0;
        pixel_data[94][190] = 0;
        pixel_data[94][191] = 0;
        pixel_data[94][192] = 0;
        pixel_data[94][193] = 0;
        pixel_data[94][194] = 0;
        pixel_data[94][195] = 0;
        pixel_data[94][196] = 0;
        pixel_data[94][197] = 0;
        pixel_data[94][198] = 0;
        pixel_data[94][199] = 0; // y=94
        pixel_data[95][0] = 0;
        pixel_data[95][1] = 0;
        pixel_data[95][2] = 0;
        pixel_data[95][3] = 0;
        pixel_data[95][4] = 0;
        pixel_data[95][5] = 0;
        pixel_data[95][6] = 0;
        pixel_data[95][7] = 0;
        pixel_data[95][8] = 0;
        pixel_data[95][9] = 0;
        pixel_data[95][10] = 0;
        pixel_data[95][11] = 0;
        pixel_data[95][12] = 0;
        pixel_data[95][13] = 0;
        pixel_data[95][14] = 0;
        pixel_data[95][15] = 0;
        pixel_data[95][16] = 0;
        pixel_data[95][17] = 0;
        pixel_data[95][18] = 0;
        pixel_data[95][19] = 0;
        pixel_data[95][20] = 0;
        pixel_data[95][21] = 0;
        pixel_data[95][22] = 0;
        pixel_data[95][23] = 0;
        pixel_data[95][24] = 0;
        pixel_data[95][25] = 0;
        pixel_data[95][26] = 0;
        pixel_data[95][27] = 0;
        pixel_data[95][28] = 0;
        pixel_data[95][29] = 0;
        pixel_data[95][30] = 0;
        pixel_data[95][31] = 0;
        pixel_data[95][32] = 0;
        pixel_data[95][33] = 0;
        pixel_data[95][34] = 0;
        pixel_data[95][35] = 0;
        pixel_data[95][36] = 0;
        pixel_data[95][37] = 0;
        pixel_data[95][38] = 0;
        pixel_data[95][39] = 0;
        pixel_data[95][40] = 0;
        pixel_data[95][41] = 0;
        pixel_data[95][42] = 0;
        pixel_data[95][43] = 0;
        pixel_data[95][44] = 0;
        pixel_data[95][45] = 0;
        pixel_data[95][46] = 0;
        pixel_data[95][47] = 0;
        pixel_data[95][48] = 0;
        pixel_data[95][49] = 0;
        pixel_data[95][50] = 0;
        pixel_data[95][51] = 0;
        pixel_data[95][52] = 0;
        pixel_data[95][53] = 0;
        pixel_data[95][54] = 0;
        pixel_data[95][55] = 0;
        pixel_data[95][56] = 0;
        pixel_data[95][57] = 0;
        pixel_data[95][58] = 0;
        pixel_data[95][59] = 0;
        pixel_data[95][60] = 0;
        pixel_data[95][61] = 0;
        pixel_data[95][62] = 0;
        pixel_data[95][63] = 0;
        pixel_data[95][64] = 0;
        pixel_data[95][65] = 0;
        pixel_data[95][66] = 0;
        pixel_data[95][67] = 0;
        pixel_data[95][68] = 0;
        pixel_data[95][69] = 0;
        pixel_data[95][70] = 0;
        pixel_data[95][71] = 0;
        pixel_data[95][72] = 0;
        pixel_data[95][73] = 0;
        pixel_data[95][74] = 0;
        pixel_data[95][75] = 0;
        pixel_data[95][76] = 0;
        pixel_data[95][77] = 0;
        pixel_data[95][78] = 0;
        pixel_data[95][79] = 0;
        pixel_data[95][80] = 0;
        pixel_data[95][81] = 0;
        pixel_data[95][82] = 0;
        pixel_data[95][83] = 0;
        pixel_data[95][84] = 0;
        pixel_data[95][85] = 0;
        pixel_data[95][86] = 0;
        pixel_data[95][87] = 0;
        pixel_data[95][88] = 0;
        pixel_data[95][89] = 0;
        pixel_data[95][90] = 0;
        pixel_data[95][91] = 0;
        pixel_data[95][92] = 0;
        pixel_data[95][93] = 0;
        pixel_data[95][94] = 0;
        pixel_data[95][95] = 0;
        pixel_data[95][96] = 0;
        pixel_data[95][97] = 0;
        pixel_data[95][98] = 0;
        pixel_data[95][99] = 0;
        pixel_data[95][100] = 0;
        pixel_data[95][101] = 0;
        pixel_data[95][102] = 0;
        pixel_data[95][103] = 0;
        pixel_data[95][104] = 0;
        pixel_data[95][105] = 0;
        pixel_data[95][106] = 0;
        pixel_data[95][107] = 0;
        pixel_data[95][108] = 0;
        pixel_data[95][109] = 0;
        pixel_data[95][110] = 0;
        pixel_data[95][111] = 0;
        pixel_data[95][112] = 0;
        pixel_data[95][113] = 0;
        pixel_data[95][114] = 0;
        pixel_data[95][115] = 0;
        pixel_data[95][116] = 0;
        pixel_data[95][117] = 0;
        pixel_data[95][118] = 0;
        pixel_data[95][119] = 0;
        pixel_data[95][120] = 0;
        pixel_data[95][121] = 0;
        pixel_data[95][122] = 0;
        pixel_data[95][123] = 0;
        pixel_data[95][124] = 0;
        pixel_data[95][125] = 0;
        pixel_data[95][126] = 0;
        pixel_data[95][127] = 0;
        pixel_data[95][128] = 0;
        pixel_data[95][129] = 0;
        pixel_data[95][130] = 0;
        pixel_data[95][131] = 0;
        pixel_data[95][132] = 0;
        pixel_data[95][133] = 0;
        pixel_data[95][134] = 0;
        pixel_data[95][135] = 0;
        pixel_data[95][136] = 0;
        pixel_data[95][137] = 0;
        pixel_data[95][138] = 0;
        pixel_data[95][139] = 0;
        pixel_data[95][140] = 0;
        pixel_data[95][141] = 0;
        pixel_data[95][142] = 0;
        pixel_data[95][143] = 0;
        pixel_data[95][144] = 0;
        pixel_data[95][145] = 0;
        pixel_data[95][146] = 0;
        pixel_data[95][147] = 0;
        pixel_data[95][148] = 0;
        pixel_data[95][149] = 0;
        pixel_data[95][150] = 0;
        pixel_data[95][151] = 0;
        pixel_data[95][152] = 0;
        pixel_data[95][153] = 0;
        pixel_data[95][154] = 0;
        pixel_data[95][155] = 0;
        pixel_data[95][156] = 0;
        pixel_data[95][157] = 0;
        pixel_data[95][158] = 0;
        pixel_data[95][159] = 0;
        pixel_data[95][160] = 0;
        pixel_data[95][161] = 0;
        pixel_data[95][162] = 0;
        pixel_data[95][163] = 0;
        pixel_data[95][164] = 0;
        pixel_data[95][165] = 0;
        pixel_data[95][166] = 0;
        pixel_data[95][167] = 0;
        pixel_data[95][168] = 0;
        pixel_data[95][169] = 0;
        pixel_data[95][170] = 0;
        pixel_data[95][171] = 0;
        pixel_data[95][172] = 0;
        pixel_data[95][173] = 0;
        pixel_data[95][174] = 0;
        pixel_data[95][175] = 0;
        pixel_data[95][176] = 0;
        pixel_data[95][177] = 0;
        pixel_data[95][178] = 0;
        pixel_data[95][179] = 0;
        pixel_data[95][180] = 0;
        pixel_data[95][181] = 0;
        pixel_data[95][182] = 0;
        pixel_data[95][183] = 0;
        pixel_data[95][184] = 0;
        pixel_data[95][185] = 0;
        pixel_data[95][186] = 0;
        pixel_data[95][187] = 0;
        pixel_data[95][188] = 0;
        pixel_data[95][189] = 0;
        pixel_data[95][190] = 0;
        pixel_data[95][191] = 0;
        pixel_data[95][192] = 0;
        pixel_data[95][193] = 0;
        pixel_data[95][194] = 0;
        pixel_data[95][195] = 0;
        pixel_data[95][196] = 0;
        pixel_data[95][197] = 0;
        pixel_data[95][198] = 0;
        pixel_data[95][199] = 0; // y=95
        pixel_data[96][0] = 0;
        pixel_data[96][1] = 0;
        pixel_data[96][2] = 0;
        pixel_data[96][3] = 0;
        pixel_data[96][4] = 0;
        pixel_data[96][5] = 0;
        pixel_data[96][6] = 0;
        pixel_data[96][7] = 0;
        pixel_data[96][8] = 0;
        pixel_data[96][9] = 0;
        pixel_data[96][10] = 0;
        pixel_data[96][11] = 0;
        pixel_data[96][12] = 0;
        pixel_data[96][13] = 0;
        pixel_data[96][14] = 0;
        pixel_data[96][15] = 0;
        pixel_data[96][16] = 0;
        pixel_data[96][17] = 0;
        pixel_data[96][18] = 0;
        pixel_data[96][19] = 0;
        pixel_data[96][20] = 0;
        pixel_data[96][21] = 0;
        pixel_data[96][22] = 0;
        pixel_data[96][23] = 0;
        pixel_data[96][24] = 0;
        pixel_data[96][25] = 0;
        pixel_data[96][26] = 0;
        pixel_data[96][27] = 0;
        pixel_data[96][28] = 0;
        pixel_data[96][29] = 0;
        pixel_data[96][30] = 0;
        pixel_data[96][31] = 0;
        pixel_data[96][32] = 0;
        pixel_data[96][33] = 0;
        pixel_data[96][34] = 0;
        pixel_data[96][35] = 0;
        pixel_data[96][36] = 0;
        pixel_data[96][37] = 0;
        pixel_data[96][38] = 0;
        pixel_data[96][39] = 0;
        pixel_data[96][40] = 0;
        pixel_data[96][41] = 0;
        pixel_data[96][42] = 0;
        pixel_data[96][43] = 0;
        pixel_data[96][44] = 0;
        pixel_data[96][45] = 0;
        pixel_data[96][46] = 0;
        pixel_data[96][47] = 0;
        pixel_data[96][48] = 0;
        pixel_data[96][49] = 0;
        pixel_data[96][50] = 0;
        pixel_data[96][51] = 0;
        pixel_data[96][52] = 0;
        pixel_data[96][53] = 0;
        pixel_data[96][54] = 0;
        pixel_data[96][55] = 0;
        pixel_data[96][56] = 0;
        pixel_data[96][57] = 0;
        pixel_data[96][58] = 0;
        pixel_data[96][59] = 0;
        pixel_data[96][60] = 0;
        pixel_data[96][61] = 0;
        pixel_data[96][62] = 0;
        pixel_data[96][63] = 0;
        pixel_data[96][64] = 0;
        pixel_data[96][65] = 0;
        pixel_data[96][66] = 0;
        pixel_data[96][67] = 0;
        pixel_data[96][68] = 0;
        pixel_data[96][69] = 0;
        pixel_data[96][70] = 0;
        pixel_data[96][71] = 0;
        pixel_data[96][72] = 0;
        pixel_data[96][73] = 0;
        pixel_data[96][74] = 0;
        pixel_data[96][75] = 0;
        pixel_data[96][76] = 0;
        pixel_data[96][77] = 0;
        pixel_data[96][78] = 0;
        pixel_data[96][79] = 0;
        pixel_data[96][80] = 0;
        pixel_data[96][81] = 0;
        pixel_data[96][82] = 0;
        pixel_data[96][83] = 0;
        pixel_data[96][84] = 0;
        pixel_data[96][85] = 0;
        pixel_data[96][86] = 0;
        pixel_data[96][87] = 0;
        pixel_data[96][88] = 0;
        pixel_data[96][89] = 0;
        pixel_data[96][90] = 0;
        pixel_data[96][91] = 0;
        pixel_data[96][92] = 0;
        pixel_data[96][93] = 0;
        pixel_data[96][94] = 0;
        pixel_data[96][95] = 0;
        pixel_data[96][96] = 0;
        pixel_data[96][97] = 0;
        pixel_data[96][98] = 0;
        pixel_data[96][99] = 0;
        pixel_data[96][100] = 0;
        pixel_data[96][101] = 0;
        pixel_data[96][102] = 0;
        pixel_data[96][103] = 0;
        pixel_data[96][104] = 0;
        pixel_data[96][105] = 0;
        pixel_data[96][106] = 0;
        pixel_data[96][107] = 0;
        pixel_data[96][108] = 0;
        pixel_data[96][109] = 0;
        pixel_data[96][110] = 0;
        pixel_data[96][111] = 0;
        pixel_data[96][112] = 0;
        pixel_data[96][113] = 0;
        pixel_data[96][114] = 0;
        pixel_data[96][115] = 0;
        pixel_data[96][116] = 0;
        pixel_data[96][117] = 0;
        pixel_data[96][118] = 0;
        pixel_data[96][119] = 0;
        pixel_data[96][120] = 0;
        pixel_data[96][121] = 0;
        pixel_data[96][122] = 0;
        pixel_data[96][123] = 0;
        pixel_data[96][124] = 0;
        pixel_data[96][125] = 0;
        pixel_data[96][126] = 0;
        pixel_data[96][127] = 0;
        pixel_data[96][128] = 0;
        pixel_data[96][129] = 0;
        pixel_data[96][130] = 0;
        pixel_data[96][131] = 0;
        pixel_data[96][132] = 0;
        pixel_data[96][133] = 0;
        pixel_data[96][134] = 0;
        pixel_data[96][135] = 0;
        pixel_data[96][136] = 0;
        pixel_data[96][137] = 0;
        pixel_data[96][138] = 0;
        pixel_data[96][139] = 0;
        pixel_data[96][140] = 0;
        pixel_data[96][141] = 0;
        pixel_data[96][142] = 0;
        pixel_data[96][143] = 0;
        pixel_data[96][144] = 0;
        pixel_data[96][145] = 0;
        pixel_data[96][146] = 0;
        pixel_data[96][147] = 0;
        pixel_data[96][148] = 0;
        pixel_data[96][149] = 0;
        pixel_data[96][150] = 0;
        pixel_data[96][151] = 0;
        pixel_data[96][152] = 0;
        pixel_data[96][153] = 0;
        pixel_data[96][154] = 0;
        pixel_data[96][155] = 0;
        pixel_data[96][156] = 0;
        pixel_data[96][157] = 0;
        pixel_data[96][158] = 0;
        pixel_data[96][159] = 0;
        pixel_data[96][160] = 0;
        pixel_data[96][161] = 0;
        pixel_data[96][162] = 0;
        pixel_data[96][163] = 0;
        pixel_data[96][164] = 0;
        pixel_data[96][165] = 0;
        pixel_data[96][166] = 0;
        pixel_data[96][167] = 0;
        pixel_data[96][168] = 0;
        pixel_data[96][169] = 0;
        pixel_data[96][170] = 0;
        pixel_data[96][171] = 0;
        pixel_data[96][172] = 0;
        pixel_data[96][173] = 0;
        pixel_data[96][174] = 0;
        pixel_data[96][175] = 0;
        pixel_data[96][176] = 0;
        pixel_data[96][177] = 0;
        pixel_data[96][178] = 0;
        pixel_data[96][179] = 0;
        pixel_data[96][180] = 0;
        pixel_data[96][181] = 0;
        pixel_data[96][182] = 0;
        pixel_data[96][183] = 0;
        pixel_data[96][184] = 0;
        pixel_data[96][185] = 0;
        pixel_data[96][186] = 0;
        pixel_data[96][187] = 0;
        pixel_data[96][188] = 0;
        pixel_data[96][189] = 0;
        pixel_data[96][190] = 0;
        pixel_data[96][191] = 0;
        pixel_data[96][192] = 0;
        pixel_data[96][193] = 0;
        pixel_data[96][194] = 0;
        pixel_data[96][195] = 0;
        pixel_data[96][196] = 0;
        pixel_data[96][197] = 0;
        pixel_data[96][198] = 0;
        pixel_data[96][199] = 0; // y=96
        pixel_data[97][0] = 0;
        pixel_data[97][1] = 0;
        pixel_data[97][2] = 0;
        pixel_data[97][3] = 0;
        pixel_data[97][4] = 0;
        pixel_data[97][5] = 0;
        pixel_data[97][6] = 0;
        pixel_data[97][7] = 0;
        pixel_data[97][8] = 0;
        pixel_data[97][9] = 0;
        pixel_data[97][10] = 0;
        pixel_data[97][11] = 0;
        pixel_data[97][12] = 0;
        pixel_data[97][13] = 0;
        pixel_data[97][14] = 0;
        pixel_data[97][15] = 0;
        pixel_data[97][16] = 0;
        pixel_data[97][17] = 0;
        pixel_data[97][18] = 0;
        pixel_data[97][19] = 0;
        pixel_data[97][20] = 0;
        pixel_data[97][21] = 0;
        pixel_data[97][22] = 0;
        pixel_data[97][23] = 0;
        pixel_data[97][24] = 0;
        pixel_data[97][25] = 0;
        pixel_data[97][26] = 0;
        pixel_data[97][27] = 0;
        pixel_data[97][28] = 0;
        pixel_data[97][29] = 0;
        pixel_data[97][30] = 0;
        pixel_data[97][31] = 0;
        pixel_data[97][32] = 0;
        pixel_data[97][33] = 0;
        pixel_data[97][34] = 0;
        pixel_data[97][35] = 0;
        pixel_data[97][36] = 0;
        pixel_data[97][37] = 0;
        pixel_data[97][38] = 0;
        pixel_data[97][39] = 0;
        pixel_data[97][40] = 0;
        pixel_data[97][41] = 0;
        pixel_data[97][42] = 0;
        pixel_data[97][43] = 0;
        pixel_data[97][44] = 0;
        pixel_data[97][45] = 0;
        pixel_data[97][46] = 0;
        pixel_data[97][47] = 0;
        pixel_data[97][48] = 0;
        pixel_data[97][49] = 0;
        pixel_data[97][50] = 0;
        pixel_data[97][51] = 0;
        pixel_data[97][52] = 0;
        pixel_data[97][53] = 0;
        pixel_data[97][54] = 0;
        pixel_data[97][55] = 0;
        pixel_data[97][56] = 0;
        pixel_data[97][57] = 0;
        pixel_data[97][58] = 0;
        pixel_data[97][59] = 0;
        pixel_data[97][60] = 0;
        pixel_data[97][61] = 0;
        pixel_data[97][62] = 0;
        pixel_data[97][63] = 0;
        pixel_data[97][64] = 0;
        pixel_data[97][65] = 0;
        pixel_data[97][66] = 0;
        pixel_data[97][67] = 0;
        pixel_data[97][68] = 0;
        pixel_data[97][69] = 0;
        pixel_data[97][70] = 0;
        pixel_data[97][71] = 0;
        pixel_data[97][72] = 0;
        pixel_data[97][73] = 0;
        pixel_data[97][74] = 0;
        pixel_data[97][75] = 0;
        pixel_data[97][76] = 0;
        pixel_data[97][77] = 0;
        pixel_data[97][78] = 0;
        pixel_data[97][79] = 0;
        pixel_data[97][80] = 0;
        pixel_data[97][81] = 0;
        pixel_data[97][82] = 0;
        pixel_data[97][83] = 0;
        pixel_data[97][84] = 0;
        pixel_data[97][85] = 0;
        pixel_data[97][86] = 0;
        pixel_data[97][87] = 0;
        pixel_data[97][88] = 0;
        pixel_data[97][89] = 0;
        pixel_data[97][90] = 0;
        pixel_data[97][91] = 0;
        pixel_data[97][92] = 0;
        pixel_data[97][93] = 0;
        pixel_data[97][94] = 0;
        pixel_data[97][95] = 0;
        pixel_data[97][96] = 0;
        pixel_data[97][97] = 0;
        pixel_data[97][98] = 0;
        pixel_data[97][99] = 0;
        pixel_data[97][100] = 0;
        pixel_data[97][101] = 0;
        pixel_data[97][102] = 0;
        pixel_data[97][103] = 0;
        pixel_data[97][104] = 0;
        pixel_data[97][105] = 0;
        pixel_data[97][106] = 0;
        pixel_data[97][107] = 0;
        pixel_data[97][108] = 0;
        pixel_data[97][109] = 0;
        pixel_data[97][110] = 0;
        pixel_data[97][111] = 0;
        pixel_data[97][112] = 0;
        pixel_data[97][113] = 0;
        pixel_data[97][114] = 0;
        pixel_data[97][115] = 0;
        pixel_data[97][116] = 0;
        pixel_data[97][117] = 0;
        pixel_data[97][118] = 0;
        pixel_data[97][119] = 0;
        pixel_data[97][120] = 0;
        pixel_data[97][121] = 0;
        pixel_data[97][122] = 0;
        pixel_data[97][123] = 0;
        pixel_data[97][124] = 0;
        pixel_data[97][125] = 0;
        pixel_data[97][126] = 0;
        pixel_data[97][127] = 0;
        pixel_data[97][128] = 0;
        pixel_data[97][129] = 0;
        pixel_data[97][130] = 0;
        pixel_data[97][131] = 0;
        pixel_data[97][132] = 0;
        pixel_data[97][133] = 0;
        pixel_data[97][134] = 0;
        pixel_data[97][135] = 0;
        pixel_data[97][136] = 0;
        pixel_data[97][137] = 0;
        pixel_data[97][138] = 0;
        pixel_data[97][139] = 0;
        pixel_data[97][140] = 0;
        pixel_data[97][141] = 0;
        pixel_data[97][142] = 0;
        pixel_data[97][143] = 0;
        pixel_data[97][144] = 0;
        pixel_data[97][145] = 0;
        pixel_data[97][146] = 0;
        pixel_data[97][147] = 0;
        pixel_data[97][148] = 0;
        pixel_data[97][149] = 0;
        pixel_data[97][150] = 0;
        pixel_data[97][151] = 0;
        pixel_data[97][152] = 0;
        pixel_data[97][153] = 0;
        pixel_data[97][154] = 0;
        pixel_data[97][155] = 0;
        pixel_data[97][156] = 0;
        pixel_data[97][157] = 0;
        pixel_data[97][158] = 0;
        pixel_data[97][159] = 0;
        pixel_data[97][160] = 0;
        pixel_data[97][161] = 0;
        pixel_data[97][162] = 0;
        pixel_data[97][163] = 0;
        pixel_data[97][164] = 0;
        pixel_data[97][165] = 0;
        pixel_data[97][166] = 0;
        pixel_data[97][167] = 0;
        pixel_data[97][168] = 0;
        pixel_data[97][169] = 0;
        pixel_data[97][170] = 0;
        pixel_data[97][171] = 0;
        pixel_data[97][172] = 0;
        pixel_data[97][173] = 0;
        pixel_data[97][174] = 0;
        pixel_data[97][175] = 0;
        pixel_data[97][176] = 0;
        pixel_data[97][177] = 0;
        pixel_data[97][178] = 0;
        pixel_data[97][179] = 0;
        pixel_data[97][180] = 0;
        pixel_data[97][181] = 0;
        pixel_data[97][182] = 0;
        pixel_data[97][183] = 0;
        pixel_data[97][184] = 0;
        pixel_data[97][185] = 0;
        pixel_data[97][186] = 0;
        pixel_data[97][187] = 0;
        pixel_data[97][188] = 0;
        pixel_data[97][189] = 0;
        pixel_data[97][190] = 0;
        pixel_data[97][191] = 0;
        pixel_data[97][192] = 0;
        pixel_data[97][193] = 0;
        pixel_data[97][194] = 0;
        pixel_data[97][195] = 0;
        pixel_data[97][196] = 0;
        pixel_data[97][197] = 0;
        pixel_data[97][198] = 0;
        pixel_data[97][199] = 0; // y=97
        pixel_data[98][0] = 0;
        pixel_data[98][1] = 0;
        pixel_data[98][2] = 0;
        pixel_data[98][3] = 0;
        pixel_data[98][4] = 0;
        pixel_data[98][5] = 0;
        pixel_data[98][6] = 0;
        pixel_data[98][7] = 0;
        pixel_data[98][8] = 0;
        pixel_data[98][9] = 0;
        pixel_data[98][10] = 0;
        pixel_data[98][11] = 0;
        pixel_data[98][12] = 0;
        pixel_data[98][13] = 0;
        pixel_data[98][14] = 0;
        pixel_data[98][15] = 0;
        pixel_data[98][16] = 0;
        pixel_data[98][17] = 0;
        pixel_data[98][18] = 0;
        pixel_data[98][19] = 0;
        pixel_data[98][20] = 0;
        pixel_data[98][21] = 0;
        pixel_data[98][22] = 0;
        pixel_data[98][23] = 0;
        pixel_data[98][24] = 0;
        pixel_data[98][25] = 0;
        pixel_data[98][26] = 0;
        pixel_data[98][27] = 0;
        pixel_data[98][28] = 0;
        pixel_data[98][29] = 0;
        pixel_data[98][30] = 0;
        pixel_data[98][31] = 0;
        pixel_data[98][32] = 0;
        pixel_data[98][33] = 0;
        pixel_data[98][34] = 0;
        pixel_data[98][35] = 0;
        pixel_data[98][36] = 0;
        pixel_data[98][37] = 0;
        pixel_data[98][38] = 0;
        pixel_data[98][39] = 0;
        pixel_data[98][40] = 0;
        pixel_data[98][41] = 0;
        pixel_data[98][42] = 0;
        pixel_data[98][43] = 0;
        pixel_data[98][44] = 0;
        pixel_data[98][45] = 0;
        pixel_data[98][46] = 0;
        pixel_data[98][47] = 0;
        pixel_data[98][48] = 0;
        pixel_data[98][49] = 0;
        pixel_data[98][50] = 0;
        pixel_data[98][51] = 0;
        pixel_data[98][52] = 0;
        pixel_data[98][53] = 0;
        pixel_data[98][54] = 0;
        pixel_data[98][55] = 0;
        pixel_data[98][56] = 0;
        pixel_data[98][57] = 0;
        pixel_data[98][58] = 0;
        pixel_data[98][59] = 0;
        pixel_data[98][60] = 0;
        pixel_data[98][61] = 0;
        pixel_data[98][62] = 0;
        pixel_data[98][63] = 0;
        pixel_data[98][64] = 0;
        pixel_data[98][65] = 0;
        pixel_data[98][66] = 0;
        pixel_data[98][67] = 0;
        pixel_data[98][68] = 0;
        pixel_data[98][69] = 0;
        pixel_data[98][70] = 0;
        pixel_data[98][71] = 0;
        pixel_data[98][72] = 0;
        pixel_data[98][73] = 0;
        pixel_data[98][74] = 0;
        pixel_data[98][75] = 0;
        pixel_data[98][76] = 0;
        pixel_data[98][77] = 0;
        pixel_data[98][78] = 0;
        pixel_data[98][79] = 0;
        pixel_data[98][80] = 0;
        pixel_data[98][81] = 0;
        pixel_data[98][82] = 0;
        pixel_data[98][83] = 0;
        pixel_data[98][84] = 0;
        pixel_data[98][85] = 0;
        pixel_data[98][86] = 0;
        pixel_data[98][87] = 0;
        pixel_data[98][88] = 0;
        pixel_data[98][89] = 0;
        pixel_data[98][90] = 0;
        pixel_data[98][91] = 0;
        pixel_data[98][92] = 0;
        pixel_data[98][93] = 0;
        pixel_data[98][94] = 0;
        pixel_data[98][95] = 0;
        pixel_data[98][96] = 0;
        pixel_data[98][97] = 0;
        pixel_data[98][98] = 0;
        pixel_data[98][99] = 0;
        pixel_data[98][100] = 0;
        pixel_data[98][101] = 0;
        pixel_data[98][102] = 0;
        pixel_data[98][103] = 0;
        pixel_data[98][104] = 0;
        pixel_data[98][105] = 0;
        pixel_data[98][106] = 0;
        pixel_data[98][107] = 0;
        pixel_data[98][108] = 0;
        pixel_data[98][109] = 0;
        pixel_data[98][110] = 0;
        pixel_data[98][111] = 0;
        pixel_data[98][112] = 0;
        pixel_data[98][113] = 0;
        pixel_data[98][114] = 0;
        pixel_data[98][115] = 0;
        pixel_data[98][116] = 0;
        pixel_data[98][117] = 0;
        pixel_data[98][118] = 0;
        pixel_data[98][119] = 0;
        pixel_data[98][120] = 0;
        pixel_data[98][121] = 0;
        pixel_data[98][122] = 0;
        pixel_data[98][123] = 0;
        pixel_data[98][124] = 0;
        pixel_data[98][125] = 0;
        pixel_data[98][126] = 0;
        pixel_data[98][127] = 0;
        pixel_data[98][128] = 0;
        pixel_data[98][129] = 0;
        pixel_data[98][130] = 0;
        pixel_data[98][131] = 0;
        pixel_data[98][132] = 0;
        pixel_data[98][133] = 0;
        pixel_data[98][134] = 0;
        pixel_data[98][135] = 0;
        pixel_data[98][136] = 0;
        pixel_data[98][137] = 0;
        pixel_data[98][138] = 0;
        pixel_data[98][139] = 0;
        pixel_data[98][140] = 0;
        pixel_data[98][141] = 0;
        pixel_data[98][142] = 0;
        pixel_data[98][143] = 0;
        pixel_data[98][144] = 0;
        pixel_data[98][145] = 0;
        pixel_data[98][146] = 0;
        pixel_data[98][147] = 0;
        pixel_data[98][148] = 0;
        pixel_data[98][149] = 0;
        pixel_data[98][150] = 0;
        pixel_data[98][151] = 0;
        pixel_data[98][152] = 0;
        pixel_data[98][153] = 0;
        pixel_data[98][154] = 0;
        pixel_data[98][155] = 0;
        pixel_data[98][156] = 0;
        pixel_data[98][157] = 0;
        pixel_data[98][158] = 0;
        pixel_data[98][159] = 0;
        pixel_data[98][160] = 0;
        pixel_data[98][161] = 0;
        pixel_data[98][162] = 0;
        pixel_data[98][163] = 0;
        pixel_data[98][164] = 0;
        pixel_data[98][165] = 0;
        pixel_data[98][166] = 0;
        pixel_data[98][167] = 0;
        pixel_data[98][168] = 0;
        pixel_data[98][169] = 0;
        pixel_data[98][170] = 0;
        pixel_data[98][171] = 0;
        pixel_data[98][172] = 0;
        pixel_data[98][173] = 0;
        pixel_data[98][174] = 0;
        pixel_data[98][175] = 0;
        pixel_data[98][176] = 0;
        pixel_data[98][177] = 0;
        pixel_data[98][178] = 0;
        pixel_data[98][179] = 0;
        pixel_data[98][180] = 0;
        pixel_data[98][181] = 0;
        pixel_data[98][182] = 0;
        pixel_data[98][183] = 0;
        pixel_data[98][184] = 0;
        pixel_data[98][185] = 0;
        pixel_data[98][186] = 0;
        pixel_data[98][187] = 0;
        pixel_data[98][188] = 0;
        pixel_data[98][189] = 0;
        pixel_data[98][190] = 0;
        pixel_data[98][191] = 0;
        pixel_data[98][192] = 0;
        pixel_data[98][193] = 0;
        pixel_data[98][194] = 0;
        pixel_data[98][195] = 0;
        pixel_data[98][196] = 0;
        pixel_data[98][197] = 0;
        pixel_data[98][198] = 0;
        pixel_data[98][199] = 0; // y=98
        pixel_data[99][0] = 0;
        pixel_data[99][1] = 0;
        pixel_data[99][2] = 0;
        pixel_data[99][3] = 0;
        pixel_data[99][4] = 0;
        pixel_data[99][5] = 0;
        pixel_data[99][6] = 0;
        pixel_data[99][7] = 0;
        pixel_data[99][8] = 0;
        pixel_data[99][9] = 0;
        pixel_data[99][10] = 0;
        pixel_data[99][11] = 0;
        pixel_data[99][12] = 0;
        pixel_data[99][13] = 0;
        pixel_data[99][14] = 0;
        pixel_data[99][15] = 0;
        pixel_data[99][16] = 0;
        pixel_data[99][17] = 0;
        pixel_data[99][18] = 0;
        pixel_data[99][19] = 0;
        pixel_data[99][20] = 0;
        pixel_data[99][21] = 0;
        pixel_data[99][22] = 0;
        pixel_data[99][23] = 0;
        pixel_data[99][24] = 0;
        pixel_data[99][25] = 0;
        pixel_data[99][26] = 0;
        pixel_data[99][27] = 0;
        pixel_data[99][28] = 0;
        pixel_data[99][29] = 0;
        pixel_data[99][30] = 0;
        pixel_data[99][31] = 0;
        pixel_data[99][32] = 0;
        pixel_data[99][33] = 0;
        pixel_data[99][34] = 0;
        pixel_data[99][35] = 0;
        pixel_data[99][36] = 0;
        pixel_data[99][37] = 0;
        pixel_data[99][38] = 0;
        pixel_data[99][39] = 0;
        pixel_data[99][40] = 0;
        pixel_data[99][41] = 0;
        pixel_data[99][42] = 0;
        pixel_data[99][43] = 0;
        pixel_data[99][44] = 0;
        pixel_data[99][45] = 0;
        pixel_data[99][46] = 0;
        pixel_data[99][47] = 0;
        pixel_data[99][48] = 0;
        pixel_data[99][49] = 0;
        pixel_data[99][50] = 0;
        pixel_data[99][51] = 0;
        pixel_data[99][52] = 0;
        pixel_data[99][53] = 0;
        pixel_data[99][54] = 0;
        pixel_data[99][55] = 0;
        pixel_data[99][56] = 0;
        pixel_data[99][57] = 0;
        pixel_data[99][58] = 0;
        pixel_data[99][59] = 0;
        pixel_data[99][60] = 0;
        pixel_data[99][61] = 0;
        pixel_data[99][62] = 0;
        pixel_data[99][63] = 0;
        pixel_data[99][64] = 0;
        pixel_data[99][65] = 0;
        pixel_data[99][66] = 0;
        pixel_data[99][67] = 0;
        pixel_data[99][68] = 0;
        pixel_data[99][69] = 0;
        pixel_data[99][70] = 0;
        pixel_data[99][71] = 0;
        pixel_data[99][72] = 0;
        pixel_data[99][73] = 0;
        pixel_data[99][74] = 0;
        pixel_data[99][75] = 0;
        pixel_data[99][76] = 0;
        pixel_data[99][77] = 0;
        pixel_data[99][78] = 0;
        pixel_data[99][79] = 0;
        pixel_data[99][80] = 0;
        pixel_data[99][81] = 0;
        pixel_data[99][82] = 0;
        pixel_data[99][83] = 0;
        pixel_data[99][84] = 0;
        pixel_data[99][85] = 0;
        pixel_data[99][86] = 0;
        pixel_data[99][87] = 0;
        pixel_data[99][88] = 0;
        pixel_data[99][89] = 0;
        pixel_data[99][90] = 0;
        pixel_data[99][91] = 0;
        pixel_data[99][92] = 0;
        pixel_data[99][93] = 0;
        pixel_data[99][94] = 0;
        pixel_data[99][95] = 0;
        pixel_data[99][96] = 0;
        pixel_data[99][97] = 0;
        pixel_data[99][98] = 0;
        pixel_data[99][99] = 0;
        pixel_data[99][100] = 0;
        pixel_data[99][101] = 0;
        pixel_data[99][102] = 0;
        pixel_data[99][103] = 0;
        pixel_data[99][104] = 0;
        pixel_data[99][105] = 0;
        pixel_data[99][106] = 0;
        pixel_data[99][107] = 0;
        pixel_data[99][108] = 0;
        pixel_data[99][109] = 0;
        pixel_data[99][110] = 0;
        pixel_data[99][111] = 0;
        pixel_data[99][112] = 0;
        pixel_data[99][113] = 0;
        pixel_data[99][114] = 0;
        pixel_data[99][115] = 0;
        pixel_data[99][116] = 0;
        pixel_data[99][117] = 0;
        pixel_data[99][118] = 0;
        pixel_data[99][119] = 0;
        pixel_data[99][120] = 0;
        pixel_data[99][121] = 0;
        pixel_data[99][122] = 0;
        pixel_data[99][123] = 0;
        pixel_data[99][124] = 0;
        pixel_data[99][125] = 0;
        pixel_data[99][126] = 0;
        pixel_data[99][127] = 0;
        pixel_data[99][128] = 0;
        pixel_data[99][129] = 0;
        pixel_data[99][130] = 0;
        pixel_data[99][131] = 0;
        pixel_data[99][132] = 0;
        pixel_data[99][133] = 0;
        pixel_data[99][134] = 0;
        pixel_data[99][135] = 0;
        pixel_data[99][136] = 0;
        pixel_data[99][137] = 0;
        pixel_data[99][138] = 0;
        pixel_data[99][139] = 0;
        pixel_data[99][140] = 0;
        pixel_data[99][141] = 0;
        pixel_data[99][142] = 0;
        pixel_data[99][143] = 0;
        pixel_data[99][144] = 0;
        pixel_data[99][145] = 0;
        pixel_data[99][146] = 0;
        pixel_data[99][147] = 0;
        pixel_data[99][148] = 0;
        pixel_data[99][149] = 0;
        pixel_data[99][150] = 0;
        pixel_data[99][151] = 0;
        pixel_data[99][152] = 0;
        pixel_data[99][153] = 0;
        pixel_data[99][154] = 0;
        pixel_data[99][155] = 0;
        pixel_data[99][156] = 0;
        pixel_data[99][157] = 0;
        pixel_data[99][158] = 0;
        pixel_data[99][159] = 0;
        pixel_data[99][160] = 0;
        pixel_data[99][161] = 0;
        pixel_data[99][162] = 0;
        pixel_data[99][163] = 0;
        pixel_data[99][164] = 0;
        pixel_data[99][165] = 0;
        pixel_data[99][166] = 0;
        pixel_data[99][167] = 0;
        pixel_data[99][168] = 0;
        pixel_data[99][169] = 0;
        pixel_data[99][170] = 0;
        pixel_data[99][171] = 0;
        pixel_data[99][172] = 0;
        pixel_data[99][173] = 0;
        pixel_data[99][174] = 0;
        pixel_data[99][175] = 0;
        pixel_data[99][176] = 0;
        pixel_data[99][177] = 0;
        pixel_data[99][178] = 0;
        pixel_data[99][179] = 0;
        pixel_data[99][180] = 0;
        pixel_data[99][181] = 0;
        pixel_data[99][182] = 0;
        pixel_data[99][183] = 0;
        pixel_data[99][184] = 0;
        pixel_data[99][185] = 0;
        pixel_data[99][186] = 0;
        pixel_data[99][187] = 0;
        pixel_data[99][188] = 0;
        pixel_data[99][189] = 0;
        pixel_data[99][190] = 0;
        pixel_data[99][191] = 0;
        pixel_data[99][192] = 0;
        pixel_data[99][193] = 0;
        pixel_data[99][194] = 0;
        pixel_data[99][195] = 0;
        pixel_data[99][196] = 0;
        pixel_data[99][197] = 0;
        pixel_data[99][198] = 0;
        pixel_data[99][199] = 0; // y=99
        pixel_data[100][0] = 0;
        pixel_data[100][1] = 0;
        pixel_data[100][2] = 0;
        pixel_data[100][3] = 0;
        pixel_data[100][4] = 0;
        pixel_data[100][5] = 0;
        pixel_data[100][6] = 0;
        pixel_data[100][7] = 0;
        pixel_data[100][8] = 0;
        pixel_data[100][9] = 0;
        pixel_data[100][10] = 0;
        pixel_data[100][11] = 0;
        pixel_data[100][12] = 0;
        pixel_data[100][13] = 0;
        pixel_data[100][14] = 0;
        pixel_data[100][15] = 0;
        pixel_data[100][16] = 0;
        pixel_data[100][17] = 0;
        pixel_data[100][18] = 0;
        pixel_data[100][19] = 0;
        pixel_data[100][20] = 0;
        pixel_data[100][21] = 0;
        pixel_data[100][22] = 0;
        pixel_data[100][23] = 0;
        pixel_data[100][24] = 0;
        pixel_data[100][25] = 0;
        pixel_data[100][26] = 0;
        pixel_data[100][27] = 0;
        pixel_data[100][28] = 0;
        pixel_data[100][29] = 0;
        pixel_data[100][30] = 0;
        pixel_data[100][31] = 0;
        pixel_data[100][32] = 0;
        pixel_data[100][33] = 0;
        pixel_data[100][34] = 0;
        pixel_data[100][35] = 0;
        pixel_data[100][36] = 0;
        pixel_data[100][37] = 0;
        pixel_data[100][38] = 0;
        pixel_data[100][39] = 0;
        pixel_data[100][40] = 0;
        pixel_data[100][41] = 0;
        pixel_data[100][42] = 0;
        pixel_data[100][43] = 0;
        pixel_data[100][44] = 0;
        pixel_data[100][45] = 0;
        pixel_data[100][46] = 0;
        pixel_data[100][47] = 0;
        pixel_data[100][48] = 0;
        pixel_data[100][49] = 0;
        pixel_data[100][50] = 0;
        pixel_data[100][51] = 0;
        pixel_data[100][52] = 0;
        pixel_data[100][53] = 0;
        pixel_data[100][54] = 0;
        pixel_data[100][55] = 0;
        pixel_data[100][56] = 0;
        pixel_data[100][57] = 0;
        pixel_data[100][58] = 0;
        pixel_data[100][59] = 0;
        pixel_data[100][60] = 0;
        pixel_data[100][61] = 0;
        pixel_data[100][62] = 0;
        pixel_data[100][63] = 0;
        pixel_data[100][64] = 0;
        pixel_data[100][65] = 0;
        pixel_data[100][66] = 0;
        pixel_data[100][67] = 0;
        pixel_data[100][68] = 0;
        pixel_data[100][69] = 0;
        pixel_data[100][70] = 0;
        pixel_data[100][71] = 0;
        pixel_data[100][72] = 0;
        pixel_data[100][73] = 0;
        pixel_data[100][74] = 0;
        pixel_data[100][75] = 0;
        pixel_data[100][76] = 0;
        pixel_data[100][77] = 0;
        pixel_data[100][78] = 0;
        pixel_data[100][79] = 0;
        pixel_data[100][80] = 0;
        pixel_data[100][81] = 0;
        pixel_data[100][82] = 0;
        pixel_data[100][83] = 0;
        pixel_data[100][84] = 0;
        pixel_data[100][85] = 0;
        pixel_data[100][86] = 0;
        pixel_data[100][87] = 0;
        pixel_data[100][88] = 0;
        pixel_data[100][89] = 0;
        pixel_data[100][90] = 0;
        pixel_data[100][91] = 0;
        pixel_data[100][92] = 0;
        pixel_data[100][93] = 0;
        pixel_data[100][94] = 0;
        pixel_data[100][95] = 0;
        pixel_data[100][96] = 0;
        pixel_data[100][97] = 0;
        pixel_data[100][98] = 0;
        pixel_data[100][99] = 0;
        pixel_data[100][100] = 0;
        pixel_data[100][101] = 0;
        pixel_data[100][102] = 0;
        pixel_data[100][103] = 0;
        pixel_data[100][104] = 0;
        pixel_data[100][105] = 0;
        pixel_data[100][106] = 0;
        pixel_data[100][107] = 0;
        pixel_data[100][108] = 0;
        pixel_data[100][109] = 0;
        pixel_data[100][110] = 0;
        pixel_data[100][111] = 0;
        pixel_data[100][112] = 0;
        pixel_data[100][113] = 0;
        pixel_data[100][114] = 0;
        pixel_data[100][115] = 0;
        pixel_data[100][116] = 0;
        pixel_data[100][117] = 0;
        pixel_data[100][118] = 0;
        pixel_data[100][119] = 0;
        pixel_data[100][120] = 0;
        pixel_data[100][121] = 0;
        pixel_data[100][122] = 0;
        pixel_data[100][123] = 0;
        pixel_data[100][124] = 0;
        pixel_data[100][125] = 0;
        pixel_data[100][126] = 0;
        pixel_data[100][127] = 0;
        pixel_data[100][128] = 0;
        pixel_data[100][129] = 0;
        pixel_data[100][130] = 0;
        pixel_data[100][131] = 0;
        pixel_data[100][132] = 0;
        pixel_data[100][133] = 0;
        pixel_data[100][134] = 0;
        pixel_data[100][135] = 0;
        pixel_data[100][136] = 0;
        pixel_data[100][137] = 0;
        pixel_data[100][138] = 0;
        pixel_data[100][139] = 0;
        pixel_data[100][140] = 0;
        pixel_data[100][141] = 0;
        pixel_data[100][142] = 0;
        pixel_data[100][143] = 0;
        pixel_data[100][144] = 0;
        pixel_data[100][145] = 0;
        pixel_data[100][146] = 0;
        pixel_data[100][147] = 0;
        pixel_data[100][148] = 0;
        pixel_data[100][149] = 0;
        pixel_data[100][150] = 0;
        pixel_data[100][151] = 0;
        pixel_data[100][152] = 0;
        pixel_data[100][153] = 0;
        pixel_data[100][154] = 0;
        pixel_data[100][155] = 0;
        pixel_data[100][156] = 0;
        pixel_data[100][157] = 0;
        pixel_data[100][158] = 0;
        pixel_data[100][159] = 0;
        pixel_data[100][160] = 0;
        pixel_data[100][161] = 0;
        pixel_data[100][162] = 0;
        pixel_data[100][163] = 0;
        pixel_data[100][164] = 0;
        pixel_data[100][165] = 0;
        pixel_data[100][166] = 0;
        pixel_data[100][167] = 0;
        pixel_data[100][168] = 0;
        pixel_data[100][169] = 0;
        pixel_data[100][170] = 0;
        pixel_data[100][171] = 0;
        pixel_data[100][172] = 0;
        pixel_data[100][173] = 0;
        pixel_data[100][174] = 0;
        pixel_data[100][175] = 0;
        pixel_data[100][176] = 0;
        pixel_data[100][177] = 0;
        pixel_data[100][178] = 0;
        pixel_data[100][179] = 0;
        pixel_data[100][180] = 0;
        pixel_data[100][181] = 0;
        pixel_data[100][182] = 0;
        pixel_data[100][183] = 0;
        pixel_data[100][184] = 0;
        pixel_data[100][185] = 0;
        pixel_data[100][186] = 0;
        pixel_data[100][187] = 0;
        pixel_data[100][188] = 0;
        pixel_data[100][189] = 0;
        pixel_data[100][190] = 0;
        pixel_data[100][191] = 0;
        pixel_data[100][192] = 0;
        pixel_data[100][193] = 0;
        pixel_data[100][194] = 0;
        pixel_data[100][195] = 0;
        pixel_data[100][196] = 0;
        pixel_data[100][197] = 0;
        pixel_data[100][198] = 0;
        pixel_data[100][199] = 0; // y=100
        pixel_data[101][0] = 0;
        pixel_data[101][1] = 0;
        pixel_data[101][2] = 0;
        pixel_data[101][3] = 0;
        pixel_data[101][4] = 0;
        pixel_data[101][5] = 0;
        pixel_data[101][6] = 0;
        pixel_data[101][7] = 0;
        pixel_data[101][8] = 0;
        pixel_data[101][9] = 0;
        pixel_data[101][10] = 0;
        pixel_data[101][11] = 0;
        pixel_data[101][12] = 0;
        pixel_data[101][13] = 0;
        pixel_data[101][14] = 0;
        pixel_data[101][15] = 0;
        pixel_data[101][16] = 0;
        pixel_data[101][17] = 0;
        pixel_data[101][18] = 0;
        pixel_data[101][19] = 0;
        pixel_data[101][20] = 0;
        pixel_data[101][21] = 0;
        pixel_data[101][22] = 0;
        pixel_data[101][23] = 0;
        pixel_data[101][24] = 0;
        pixel_data[101][25] = 0;
        pixel_data[101][26] = 0;
        pixel_data[101][27] = 0;
        pixel_data[101][28] = 0;
        pixel_data[101][29] = 0;
        pixel_data[101][30] = 0;
        pixel_data[101][31] = 0;
        pixel_data[101][32] = 0;
        pixel_data[101][33] = 0;
        pixel_data[101][34] = 0;
        pixel_data[101][35] = 0;
        pixel_data[101][36] = 0;
        pixel_data[101][37] = 0;
        pixel_data[101][38] = 0;
        pixel_data[101][39] = 0;
        pixel_data[101][40] = 0;
        pixel_data[101][41] = 0;
        pixel_data[101][42] = 0;
        pixel_data[101][43] = 0;
        pixel_data[101][44] = 0;
        pixel_data[101][45] = 0;
        pixel_data[101][46] = 0;
        pixel_data[101][47] = 0;
        pixel_data[101][48] = 0;
        pixel_data[101][49] = 0;
        pixel_data[101][50] = 0;
        pixel_data[101][51] = 0;
        pixel_data[101][52] = 0;
        pixel_data[101][53] = 0;
        pixel_data[101][54] = 0;
        pixel_data[101][55] = 0;
        pixel_data[101][56] = 0;
        pixel_data[101][57] = 0;
        pixel_data[101][58] = 0;
        pixel_data[101][59] = 0;
        pixel_data[101][60] = 0;
        pixel_data[101][61] = 0;
        pixel_data[101][62] = 0;
        pixel_data[101][63] = 0;
        pixel_data[101][64] = 0;
        pixel_data[101][65] = 0;
        pixel_data[101][66] = 0;
        pixel_data[101][67] = 0;
        pixel_data[101][68] = 0;
        pixel_data[101][69] = 0;
        pixel_data[101][70] = 0;
        pixel_data[101][71] = 0;
        pixel_data[101][72] = 0;
        pixel_data[101][73] = 0;
        pixel_data[101][74] = 0;
        pixel_data[101][75] = 0;
        pixel_data[101][76] = 0;
        pixel_data[101][77] = 0;
        pixel_data[101][78] = 0;
        pixel_data[101][79] = 0;
        pixel_data[101][80] = 0;
        pixel_data[101][81] = 0;
        pixel_data[101][82] = 0;
        pixel_data[101][83] = 0;
        pixel_data[101][84] = 0;
        pixel_data[101][85] = 0;
        pixel_data[101][86] = 0;
        pixel_data[101][87] = 0;
        pixel_data[101][88] = 0;
        pixel_data[101][89] = 0;
        pixel_data[101][90] = 0;
        pixel_data[101][91] = 0;
        pixel_data[101][92] = 0;
        pixel_data[101][93] = 0;
        pixel_data[101][94] = 0;
        pixel_data[101][95] = 0;
        pixel_data[101][96] = 0;
        pixel_data[101][97] = 0;
        pixel_data[101][98] = 0;
        pixel_data[101][99] = 0;
        pixel_data[101][100] = 0;
        pixel_data[101][101] = 0;
        pixel_data[101][102] = 0;
        pixel_data[101][103] = 0;
        pixel_data[101][104] = 0;
        pixel_data[101][105] = 0;
        pixel_data[101][106] = 0;
        pixel_data[101][107] = 0;
        pixel_data[101][108] = 0;
        pixel_data[101][109] = 0;
        pixel_data[101][110] = 0;
        pixel_data[101][111] = 0;
        pixel_data[101][112] = 0;
        pixel_data[101][113] = 0;
        pixel_data[101][114] = 0;
        pixel_data[101][115] = 0;
        pixel_data[101][116] = 0;
        pixel_data[101][117] = 0;
        pixel_data[101][118] = 0;
        pixel_data[101][119] = 0;
        pixel_data[101][120] = 0;
        pixel_data[101][121] = 0;
        pixel_data[101][122] = 0;
        pixel_data[101][123] = 0;
        pixel_data[101][124] = 0;
        pixel_data[101][125] = 0;
        pixel_data[101][126] = 0;
        pixel_data[101][127] = 0;
        pixel_data[101][128] = 0;
        pixel_data[101][129] = 0;
        pixel_data[101][130] = 0;
        pixel_data[101][131] = 0;
        pixel_data[101][132] = 0;
        pixel_data[101][133] = 0;
        pixel_data[101][134] = 0;
        pixel_data[101][135] = 0;
        pixel_data[101][136] = 0;
        pixel_data[101][137] = 0;
        pixel_data[101][138] = 0;
        pixel_data[101][139] = 0;
        pixel_data[101][140] = 0;
        pixel_data[101][141] = 0;
        pixel_data[101][142] = 0;
        pixel_data[101][143] = 0;
        pixel_data[101][144] = 0;
        pixel_data[101][145] = 0;
        pixel_data[101][146] = 0;
        pixel_data[101][147] = 0;
        pixel_data[101][148] = 0;
        pixel_data[101][149] = 0;
        pixel_data[101][150] = 0;
        pixel_data[101][151] = 0;
        pixel_data[101][152] = 0;
        pixel_data[101][153] = 0;
        pixel_data[101][154] = 0;
        pixel_data[101][155] = 0;
        pixel_data[101][156] = 0;
        pixel_data[101][157] = 0;
        pixel_data[101][158] = 0;
        pixel_data[101][159] = 0;
        pixel_data[101][160] = 0;
        pixel_data[101][161] = 0;
        pixel_data[101][162] = 0;
        pixel_data[101][163] = 0;
        pixel_data[101][164] = 0;
        pixel_data[101][165] = 0;
        pixel_data[101][166] = 0;
        pixel_data[101][167] = 0;
        pixel_data[101][168] = 0;
        pixel_data[101][169] = 0;
        pixel_data[101][170] = 0;
        pixel_data[101][171] = 0;
        pixel_data[101][172] = 0;
        pixel_data[101][173] = 0;
        pixel_data[101][174] = 0;
        pixel_data[101][175] = 0;
        pixel_data[101][176] = 0;
        pixel_data[101][177] = 0;
        pixel_data[101][178] = 0;
        pixel_data[101][179] = 0;
        pixel_data[101][180] = 0;
        pixel_data[101][181] = 0;
        pixel_data[101][182] = 0;
        pixel_data[101][183] = 0;
        pixel_data[101][184] = 0;
        pixel_data[101][185] = 0;
        pixel_data[101][186] = 0;
        pixel_data[101][187] = 0;
        pixel_data[101][188] = 0;
        pixel_data[101][189] = 0;
        pixel_data[101][190] = 0;
        pixel_data[101][191] = 0;
        pixel_data[101][192] = 0;
        pixel_data[101][193] = 0;
        pixel_data[101][194] = 0;
        pixel_data[101][195] = 0;
        pixel_data[101][196] = 0;
        pixel_data[101][197] = 0;
        pixel_data[101][198] = 0;
        pixel_data[101][199] = 0; // y=101
        pixel_data[102][0] = 0;
        pixel_data[102][1] = 0;
        pixel_data[102][2] = 0;
        pixel_data[102][3] = 0;
        pixel_data[102][4] = 0;
        pixel_data[102][5] = 0;
        pixel_data[102][6] = 0;
        pixel_data[102][7] = 0;
        pixel_data[102][8] = 0;
        pixel_data[102][9] = 0;
        pixel_data[102][10] = 0;
        pixel_data[102][11] = 0;
        pixel_data[102][12] = 0;
        pixel_data[102][13] = 0;
        pixel_data[102][14] = 0;
        pixel_data[102][15] = 0;
        pixel_data[102][16] = 0;
        pixel_data[102][17] = 0;
        pixel_data[102][18] = 0;
        pixel_data[102][19] = 0;
        pixel_data[102][20] = 0;
        pixel_data[102][21] = 0;
        pixel_data[102][22] = 0;
        pixel_data[102][23] = 0;
        pixel_data[102][24] = 0;
        pixel_data[102][25] = 0;
        pixel_data[102][26] = 0;
        pixel_data[102][27] = 0;
        pixel_data[102][28] = 0;
        pixel_data[102][29] = 0;
        pixel_data[102][30] = 0;
        pixel_data[102][31] = 0;
        pixel_data[102][32] = 0;
        pixel_data[102][33] = 0;
        pixel_data[102][34] = 0;
        pixel_data[102][35] = 0;
        pixel_data[102][36] = 0;
        pixel_data[102][37] = 0;
        pixel_data[102][38] = 0;
        pixel_data[102][39] = 0;
        pixel_data[102][40] = 0;
        pixel_data[102][41] = 0;
        pixel_data[102][42] = 0;
        pixel_data[102][43] = 0;
        pixel_data[102][44] = 0;
        pixel_data[102][45] = 0;
        pixel_data[102][46] = 0;
        pixel_data[102][47] = 0;
        pixel_data[102][48] = 0;
        pixel_data[102][49] = 0;
        pixel_data[102][50] = 0;
        pixel_data[102][51] = 0;
        pixel_data[102][52] = 0;
        pixel_data[102][53] = 0;
        pixel_data[102][54] = 0;
        pixel_data[102][55] = 0;
        pixel_data[102][56] = 0;
        pixel_data[102][57] = 0;
        pixel_data[102][58] = 0;
        pixel_data[102][59] = 0;
        pixel_data[102][60] = 0;
        pixel_data[102][61] = 0;
        pixel_data[102][62] = 0;
        pixel_data[102][63] = 0;
        pixel_data[102][64] = 0;
        pixel_data[102][65] = 0;
        pixel_data[102][66] = 0;
        pixel_data[102][67] = 0;
        pixel_data[102][68] = 0;
        pixel_data[102][69] = 0;
        pixel_data[102][70] = 0;
        pixel_data[102][71] = 0;
        pixel_data[102][72] = 0;
        pixel_data[102][73] = 0;
        pixel_data[102][74] = 0;
        pixel_data[102][75] = 0;
        pixel_data[102][76] = 0;
        pixel_data[102][77] = 0;
        pixel_data[102][78] = 0;
        pixel_data[102][79] = 0;
        pixel_data[102][80] = 0;
        pixel_data[102][81] = 0;
        pixel_data[102][82] = 0;
        pixel_data[102][83] = 0;
        pixel_data[102][84] = 0;
        pixel_data[102][85] = 0;
        pixel_data[102][86] = 0;
        pixel_data[102][87] = 0;
        pixel_data[102][88] = 0;
        pixel_data[102][89] = 0;
        pixel_data[102][90] = 0;
        pixel_data[102][91] = 0;
        pixel_data[102][92] = 0;
        pixel_data[102][93] = 0;
        pixel_data[102][94] = 0;
        pixel_data[102][95] = 0;
        pixel_data[102][96] = 0;
        pixel_data[102][97] = 0;
        pixel_data[102][98] = 0;
        pixel_data[102][99] = 0;
        pixel_data[102][100] = 0;
        pixel_data[102][101] = 0;
        pixel_data[102][102] = 0;
        pixel_data[102][103] = 0;
        pixel_data[102][104] = 0;
        pixel_data[102][105] = 0;
        pixel_data[102][106] = 0;
        pixel_data[102][107] = 0;
        pixel_data[102][108] = 0;
        pixel_data[102][109] = 0;
        pixel_data[102][110] = 0;
        pixel_data[102][111] = 0;
        pixel_data[102][112] = 0;
        pixel_data[102][113] = 0;
        pixel_data[102][114] = 0;
        pixel_data[102][115] = 0;
        pixel_data[102][116] = 0;
        pixel_data[102][117] = 0;
        pixel_data[102][118] = 0;
        pixel_data[102][119] = 0;
        pixel_data[102][120] = 0;
        pixel_data[102][121] = 0;
        pixel_data[102][122] = 0;
        pixel_data[102][123] = 0;
        pixel_data[102][124] = 0;
        pixel_data[102][125] = 0;
        pixel_data[102][126] = 0;
        pixel_data[102][127] = 0;
        pixel_data[102][128] = 0;
        pixel_data[102][129] = 0;
        pixel_data[102][130] = 0;
        pixel_data[102][131] = 0;
        pixel_data[102][132] = 0;
        pixel_data[102][133] = 0;
        pixel_data[102][134] = 0;
        pixel_data[102][135] = 0;
        pixel_data[102][136] = 0;
        pixel_data[102][137] = 0;
        pixel_data[102][138] = 0;
        pixel_data[102][139] = 0;
        pixel_data[102][140] = 0;
        pixel_data[102][141] = 0;
        pixel_data[102][142] = 0;
        pixel_data[102][143] = 0;
        pixel_data[102][144] = 0;
        pixel_data[102][145] = 0;
        pixel_data[102][146] = 0;
        pixel_data[102][147] = 0;
        pixel_data[102][148] = 0;
        pixel_data[102][149] = 0;
        pixel_data[102][150] = 0;
        pixel_data[102][151] = 0;
        pixel_data[102][152] = 0;
        pixel_data[102][153] = 0;
        pixel_data[102][154] = 0;
        pixel_data[102][155] = 0;
        pixel_data[102][156] = 0;
        pixel_data[102][157] = 0;
        pixel_data[102][158] = 0;
        pixel_data[102][159] = 0;
        pixel_data[102][160] = 0;
        pixel_data[102][161] = 0;
        pixel_data[102][162] = 0;
        pixel_data[102][163] = 0;
        pixel_data[102][164] = 0;
        pixel_data[102][165] = 0;
        pixel_data[102][166] = 0;
        pixel_data[102][167] = 0;
        pixel_data[102][168] = 0;
        pixel_data[102][169] = 0;
        pixel_data[102][170] = 0;
        pixel_data[102][171] = 0;
        pixel_data[102][172] = 0;
        pixel_data[102][173] = 0;
        pixel_data[102][174] = 0;
        pixel_data[102][175] = 0;
        pixel_data[102][176] = 0;
        pixel_data[102][177] = 0;
        pixel_data[102][178] = 0;
        pixel_data[102][179] = 0;
        pixel_data[102][180] = 0;
        pixel_data[102][181] = 0;
        pixel_data[102][182] = 0;
        pixel_data[102][183] = 0;
        pixel_data[102][184] = 0;
        pixel_data[102][185] = 0;
        pixel_data[102][186] = 0;
        pixel_data[102][187] = 0;
        pixel_data[102][188] = 0;
        pixel_data[102][189] = 0;
        pixel_data[102][190] = 0;
        pixel_data[102][191] = 0;
        pixel_data[102][192] = 0;
        pixel_data[102][193] = 0;
        pixel_data[102][194] = 0;
        pixel_data[102][195] = 0;
        pixel_data[102][196] = 0;
        pixel_data[102][197] = 0;
        pixel_data[102][198] = 0;
        pixel_data[102][199] = 0; // y=102
        pixel_data[103][0] = 0;
        pixel_data[103][1] = 0;
        pixel_data[103][2] = 0;
        pixel_data[103][3] = 0;
        pixel_data[103][4] = 0;
        pixel_data[103][5] = 0;
        pixel_data[103][6] = 0;
        pixel_data[103][7] = 0;
        pixel_data[103][8] = 0;
        pixel_data[103][9] = 0;
        pixel_data[103][10] = 0;
        pixel_data[103][11] = 0;
        pixel_data[103][12] = 0;
        pixel_data[103][13] = 0;
        pixel_data[103][14] = 0;
        pixel_data[103][15] = 0;
        pixel_data[103][16] = 0;
        pixel_data[103][17] = 0;
        pixel_data[103][18] = 0;
        pixel_data[103][19] = 0;
        pixel_data[103][20] = 0;
        pixel_data[103][21] = 0;
        pixel_data[103][22] = 0;
        pixel_data[103][23] = 0;
        pixel_data[103][24] = 0;
        pixel_data[103][25] = 0;
        pixel_data[103][26] = 0;
        pixel_data[103][27] = 0;
        pixel_data[103][28] = 0;
        pixel_data[103][29] = 0;
        pixel_data[103][30] = 0;
        pixel_data[103][31] = 0;
        pixel_data[103][32] = 0;
        pixel_data[103][33] = 0;
        pixel_data[103][34] = 0;
        pixel_data[103][35] = 0;
        pixel_data[103][36] = 0;
        pixel_data[103][37] = 0;
        pixel_data[103][38] = 0;
        pixel_data[103][39] = 0;
        pixel_data[103][40] = 0;
        pixel_data[103][41] = 0;
        pixel_data[103][42] = 0;
        pixel_data[103][43] = 0;
        pixel_data[103][44] = 0;
        pixel_data[103][45] = 0;
        pixel_data[103][46] = 0;
        pixel_data[103][47] = 0;
        pixel_data[103][48] = 0;
        pixel_data[103][49] = 0;
        pixel_data[103][50] = 0;
        pixel_data[103][51] = 0;
        pixel_data[103][52] = 0;
        pixel_data[103][53] = 0;
        pixel_data[103][54] = 0;
        pixel_data[103][55] = 0;
        pixel_data[103][56] = 0;
        pixel_data[103][57] = 0;
        pixel_data[103][58] = 0;
        pixel_data[103][59] = 0;
        pixel_data[103][60] = 0;
        pixel_data[103][61] = 0;
        pixel_data[103][62] = 0;
        pixel_data[103][63] = 0;
        pixel_data[103][64] = 0;
        pixel_data[103][65] = 0;
        pixel_data[103][66] = 0;
        pixel_data[103][67] = 0;
        pixel_data[103][68] = 0;
        pixel_data[103][69] = 0;
        pixel_data[103][70] = 0;
        pixel_data[103][71] = 0;
        pixel_data[103][72] = 0;
        pixel_data[103][73] = 0;
        pixel_data[103][74] = 0;
        pixel_data[103][75] = 0;
        pixel_data[103][76] = 0;
        pixel_data[103][77] = 0;
        pixel_data[103][78] = 0;
        pixel_data[103][79] = 0;
        pixel_data[103][80] = 0;
        pixel_data[103][81] = 0;
        pixel_data[103][82] = 0;
        pixel_data[103][83] = 0;
        pixel_data[103][84] = 0;
        pixel_data[103][85] = 0;
        pixel_data[103][86] = 0;
        pixel_data[103][87] = 0;
        pixel_data[103][88] = 0;
        pixel_data[103][89] = 0;
        pixel_data[103][90] = 0;
        pixel_data[103][91] = 0;
        pixel_data[103][92] = 0;
        pixel_data[103][93] = 0;
        pixel_data[103][94] = 0;
        pixel_data[103][95] = 0;
        pixel_data[103][96] = 0;
        pixel_data[103][97] = 0;
        pixel_data[103][98] = 0;
        pixel_data[103][99] = 0;
        pixel_data[103][100] = 0;
        pixel_data[103][101] = 0;
        pixel_data[103][102] = 0;
        pixel_data[103][103] = 0;
        pixel_data[103][104] = 0;
        pixel_data[103][105] = 0;
        pixel_data[103][106] = 0;
        pixel_data[103][107] = 0;
        pixel_data[103][108] = 0;
        pixel_data[103][109] = 0;
        pixel_data[103][110] = 0;
        pixel_data[103][111] = 0;
        pixel_data[103][112] = 0;
        pixel_data[103][113] = 0;
        pixel_data[103][114] = 0;
        pixel_data[103][115] = 0;
        pixel_data[103][116] = 0;
        pixel_data[103][117] = 0;
        pixel_data[103][118] = 0;
        pixel_data[103][119] = 0;
        pixel_data[103][120] = 0;
        pixel_data[103][121] = 0;
        pixel_data[103][122] = 0;
        pixel_data[103][123] = 0;
        pixel_data[103][124] = 0;
        pixel_data[103][125] = 0;
        pixel_data[103][126] = 0;
        pixel_data[103][127] = 0;
        pixel_data[103][128] = 0;
        pixel_data[103][129] = 0;
        pixel_data[103][130] = 0;
        pixel_data[103][131] = 0;
        pixel_data[103][132] = 0;
        pixel_data[103][133] = 0;
        pixel_data[103][134] = 0;
        pixel_data[103][135] = 0;
        pixel_data[103][136] = 0;
        pixel_data[103][137] = 0;
        pixel_data[103][138] = 0;
        pixel_data[103][139] = 0;
        pixel_data[103][140] = 0;
        pixel_data[103][141] = 0;
        pixel_data[103][142] = 0;
        pixel_data[103][143] = 0;
        pixel_data[103][144] = 0;
        pixel_data[103][145] = 0;
        pixel_data[103][146] = 0;
        pixel_data[103][147] = 0;
        pixel_data[103][148] = 0;
        pixel_data[103][149] = 0;
        pixel_data[103][150] = 0;
        pixel_data[103][151] = 0;
        pixel_data[103][152] = 0;
        pixel_data[103][153] = 0;
        pixel_data[103][154] = 0;
        pixel_data[103][155] = 0;
        pixel_data[103][156] = 0;
        pixel_data[103][157] = 0;
        pixel_data[103][158] = 0;
        pixel_data[103][159] = 0;
        pixel_data[103][160] = 0;
        pixel_data[103][161] = 0;
        pixel_data[103][162] = 0;
        pixel_data[103][163] = 0;
        pixel_data[103][164] = 0;
        pixel_data[103][165] = 0;
        pixel_data[103][166] = 0;
        pixel_data[103][167] = 0;
        pixel_data[103][168] = 0;
        pixel_data[103][169] = 0;
        pixel_data[103][170] = 0;
        pixel_data[103][171] = 0;
        pixel_data[103][172] = 0;
        pixel_data[103][173] = 0;
        pixel_data[103][174] = 0;
        pixel_data[103][175] = 0;
        pixel_data[103][176] = 0;
        pixel_data[103][177] = 0;
        pixel_data[103][178] = 0;
        pixel_data[103][179] = 0;
        pixel_data[103][180] = 0;
        pixel_data[103][181] = 0;
        pixel_data[103][182] = 0;
        pixel_data[103][183] = 0;
        pixel_data[103][184] = 0;
        pixel_data[103][185] = 0;
        pixel_data[103][186] = 0;
        pixel_data[103][187] = 0;
        pixel_data[103][188] = 0;
        pixel_data[103][189] = 0;
        pixel_data[103][190] = 0;
        pixel_data[103][191] = 0;
        pixel_data[103][192] = 0;
        pixel_data[103][193] = 0;
        pixel_data[103][194] = 0;
        pixel_data[103][195] = 0;
        pixel_data[103][196] = 0;
        pixel_data[103][197] = 0;
        pixel_data[103][198] = 0;
        pixel_data[103][199] = 0; // y=103
        pixel_data[104][0] = 0;
        pixel_data[104][1] = 0;
        pixel_data[104][2] = 0;
        pixel_data[104][3] = 0;
        pixel_data[104][4] = 0;
        pixel_data[104][5] = 0;
        pixel_data[104][6] = 0;
        pixel_data[104][7] = 0;
        pixel_data[104][8] = 0;
        pixel_data[104][9] = 0;
        pixel_data[104][10] = 0;
        pixel_data[104][11] = 0;
        pixel_data[104][12] = 0;
        pixel_data[104][13] = 0;
        pixel_data[104][14] = 0;
        pixel_data[104][15] = 0;
        pixel_data[104][16] = 0;
        pixel_data[104][17] = 0;
        pixel_data[104][18] = 0;
        pixel_data[104][19] = 0;
        pixel_data[104][20] = 0;
        pixel_data[104][21] = 0;
        pixel_data[104][22] = 0;
        pixel_data[104][23] = 0;
        pixel_data[104][24] = 0;
        pixel_data[104][25] = 0;
        pixel_data[104][26] = 0;
        pixel_data[104][27] = 0;
        pixel_data[104][28] = 0;
        pixel_data[104][29] = 0;
        pixel_data[104][30] = 0;
        pixel_data[104][31] = 0;
        pixel_data[104][32] = 0;
        pixel_data[104][33] = 0;
        pixel_data[104][34] = 0;
        pixel_data[104][35] = 0;
        pixel_data[104][36] = 0;
        pixel_data[104][37] = 0;
        pixel_data[104][38] = 0;
        pixel_data[104][39] = 0;
        pixel_data[104][40] = 0;
        pixel_data[104][41] = 0;
        pixel_data[104][42] = 0;
        pixel_data[104][43] = 0;
        pixel_data[104][44] = 0;
        pixel_data[104][45] = 0;
        pixel_data[104][46] = 0;
        pixel_data[104][47] = 0;
        pixel_data[104][48] = 0;
        pixel_data[104][49] = 0;
        pixel_data[104][50] = 0;
        pixel_data[104][51] = 0;
        pixel_data[104][52] = 0;
        pixel_data[104][53] = 0;
        pixel_data[104][54] = 0;
        pixel_data[104][55] = 0;
        pixel_data[104][56] = 0;
        pixel_data[104][57] = 0;
        pixel_data[104][58] = 0;
        pixel_data[104][59] = 0;
        pixel_data[104][60] = 0;
        pixel_data[104][61] = 0;
        pixel_data[104][62] = 0;
        pixel_data[104][63] = 0;
        pixel_data[104][64] = 0;
        pixel_data[104][65] = 0;
        pixel_data[104][66] = 0;
        pixel_data[104][67] = 0;
        pixel_data[104][68] = 0;
        pixel_data[104][69] = 0;
        pixel_data[104][70] = 0;
        pixel_data[104][71] = 0;
        pixel_data[104][72] = 0;
        pixel_data[104][73] = 0;
        pixel_data[104][74] = 0;
        pixel_data[104][75] = 0;
        pixel_data[104][76] = 0;
        pixel_data[104][77] = 0;
        pixel_data[104][78] = 0;
        pixel_data[104][79] = 0;
        pixel_data[104][80] = 0;
        pixel_data[104][81] = 0;
        pixel_data[104][82] = 0;
        pixel_data[104][83] = 0;
        pixel_data[104][84] = 0;
        pixel_data[104][85] = 0;
        pixel_data[104][86] = 0;
        pixel_data[104][87] = 0;
        pixel_data[104][88] = 0;
        pixel_data[104][89] = 0;
        pixel_data[104][90] = 0;
        pixel_data[104][91] = 0;
        pixel_data[104][92] = 0;
        pixel_data[104][93] = 0;
        pixel_data[104][94] = 0;
        pixel_data[104][95] = 0;
        pixel_data[104][96] = 0;
        pixel_data[104][97] = 0;
        pixel_data[104][98] = 0;
        pixel_data[104][99] = 0;
        pixel_data[104][100] = 0;
        pixel_data[104][101] = 0;
        pixel_data[104][102] = 0;
        pixel_data[104][103] = 0;
        pixel_data[104][104] = 0;
        pixel_data[104][105] = 0;
        pixel_data[104][106] = 0;
        pixel_data[104][107] = 0;
        pixel_data[104][108] = 0;
        pixel_data[104][109] = 0;
        pixel_data[104][110] = 0;
        pixel_data[104][111] = 0;
        pixel_data[104][112] = 0;
        pixel_data[104][113] = 0;
        pixel_data[104][114] = 0;
        pixel_data[104][115] = 0;
        pixel_data[104][116] = 0;
        pixel_data[104][117] = 0;
        pixel_data[104][118] = 0;
        pixel_data[104][119] = 0;
        pixel_data[104][120] = 0;
        pixel_data[104][121] = 0;
        pixel_data[104][122] = 0;
        pixel_data[104][123] = 0;
        pixel_data[104][124] = 0;
        pixel_data[104][125] = 0;
        pixel_data[104][126] = 0;
        pixel_data[104][127] = 0;
        pixel_data[104][128] = 0;
        pixel_data[104][129] = 0;
        pixel_data[104][130] = 0;
        pixel_data[104][131] = 0;
        pixel_data[104][132] = 0;
        pixel_data[104][133] = 0;
        pixel_data[104][134] = 0;
        pixel_data[104][135] = 0;
        pixel_data[104][136] = 0;
        pixel_data[104][137] = 0;
        pixel_data[104][138] = 0;
        pixel_data[104][139] = 0;
        pixel_data[104][140] = 0;
        pixel_data[104][141] = 0;
        pixel_data[104][142] = 0;
        pixel_data[104][143] = 0;
        pixel_data[104][144] = 0;
        pixel_data[104][145] = 0;
        pixel_data[104][146] = 0;
        pixel_data[104][147] = 0;
        pixel_data[104][148] = 0;
        pixel_data[104][149] = 0;
        pixel_data[104][150] = 0;
        pixel_data[104][151] = 0;
        pixel_data[104][152] = 0;
        pixel_data[104][153] = 0;
        pixel_data[104][154] = 0;
        pixel_data[104][155] = 0;
        pixel_data[104][156] = 0;
        pixel_data[104][157] = 0;
        pixel_data[104][158] = 0;
        pixel_data[104][159] = 0;
        pixel_data[104][160] = 0;
        pixel_data[104][161] = 0;
        pixel_data[104][162] = 0;
        pixel_data[104][163] = 0;
        pixel_data[104][164] = 0;
        pixel_data[104][165] = 0;
        pixel_data[104][166] = 0;
        pixel_data[104][167] = 0;
        pixel_data[104][168] = 0;
        pixel_data[104][169] = 0;
        pixel_data[104][170] = 0;
        pixel_data[104][171] = 0;
        pixel_data[104][172] = 0;
        pixel_data[104][173] = 0;
        pixel_data[104][174] = 0;
        pixel_data[104][175] = 0;
        pixel_data[104][176] = 0;
        pixel_data[104][177] = 0;
        pixel_data[104][178] = 0;
        pixel_data[104][179] = 0;
        pixel_data[104][180] = 0;
        pixel_data[104][181] = 0;
        pixel_data[104][182] = 0;
        pixel_data[104][183] = 0;
        pixel_data[104][184] = 0;
        pixel_data[104][185] = 0;
        pixel_data[104][186] = 0;
        pixel_data[104][187] = 0;
        pixel_data[104][188] = 0;
        pixel_data[104][189] = 0;
        pixel_data[104][190] = 0;
        pixel_data[104][191] = 0;
        pixel_data[104][192] = 0;
        pixel_data[104][193] = 0;
        pixel_data[104][194] = 0;
        pixel_data[104][195] = 0;
        pixel_data[104][196] = 0;
        pixel_data[104][197] = 0;
        pixel_data[104][198] = 0;
        pixel_data[104][199] = 0; // y=104
        pixel_data[105][0] = 0;
        pixel_data[105][1] = 0;
        pixel_data[105][2] = 0;
        pixel_data[105][3] = 0;
        pixel_data[105][4] = 0;
        pixel_data[105][5] = 0;
        pixel_data[105][6] = 0;
        pixel_data[105][7] = 0;
        pixel_data[105][8] = 0;
        pixel_data[105][9] = 0;
        pixel_data[105][10] = 0;
        pixel_data[105][11] = 0;
        pixel_data[105][12] = 0;
        pixel_data[105][13] = 0;
        pixel_data[105][14] = 0;
        pixel_data[105][15] = 0;
        pixel_data[105][16] = 0;
        pixel_data[105][17] = 0;
        pixel_data[105][18] = 0;
        pixel_data[105][19] = 0;
        pixel_data[105][20] = 0;
        pixel_data[105][21] = 0;
        pixel_data[105][22] = 0;
        pixel_data[105][23] = 0;
        pixel_data[105][24] = 0;
        pixel_data[105][25] = 0;
        pixel_data[105][26] = 0;
        pixel_data[105][27] = 0;
        pixel_data[105][28] = 0;
        pixel_data[105][29] = 0;
        pixel_data[105][30] = 0;
        pixel_data[105][31] = 0;
        pixel_data[105][32] = 0;
        pixel_data[105][33] = 0;
        pixel_data[105][34] = 0;
        pixel_data[105][35] = 0;
        pixel_data[105][36] = 0;
        pixel_data[105][37] = 0;
        pixel_data[105][38] = 0;
        pixel_data[105][39] = 0;
        pixel_data[105][40] = 0;
        pixel_data[105][41] = 0;
        pixel_data[105][42] = 0;
        pixel_data[105][43] = 0;
        pixel_data[105][44] = 0;
        pixel_data[105][45] = 0;
        pixel_data[105][46] = 0;
        pixel_data[105][47] = 0;
        pixel_data[105][48] = 0;
        pixel_data[105][49] = 0;
        pixel_data[105][50] = 0;
        pixel_data[105][51] = 0;
        pixel_data[105][52] = 0;
        pixel_data[105][53] = 0;
        pixel_data[105][54] = 0;
        pixel_data[105][55] = 0;
        pixel_data[105][56] = 0;
        pixel_data[105][57] = 0;
        pixel_data[105][58] = 0;
        pixel_data[105][59] = 0;
        pixel_data[105][60] = 0;
        pixel_data[105][61] = 0;
        pixel_data[105][62] = 0;
        pixel_data[105][63] = 0;
        pixel_data[105][64] = 0;
        pixel_data[105][65] = 0;
        pixel_data[105][66] = 0;
        pixel_data[105][67] = 0;
        pixel_data[105][68] = 0;
        pixel_data[105][69] = 0;
        pixel_data[105][70] = 0;
        pixel_data[105][71] = 0;
        pixel_data[105][72] = 0;
        pixel_data[105][73] = 0;
        pixel_data[105][74] = 0;
        pixel_data[105][75] = 0;
        pixel_data[105][76] = 0;
        pixel_data[105][77] = 0;
        pixel_data[105][78] = 0;
        pixel_data[105][79] = 0;
        pixel_data[105][80] = 0;
        pixel_data[105][81] = 0;
        pixel_data[105][82] = 0;
        pixel_data[105][83] = 0;
        pixel_data[105][84] = 0;
        pixel_data[105][85] = 0;
        pixel_data[105][86] = 0;
        pixel_data[105][87] = 0;
        pixel_data[105][88] = 0;
        pixel_data[105][89] = 0;
        pixel_data[105][90] = 0;
        pixel_data[105][91] = 0;
        pixel_data[105][92] = 0;
        pixel_data[105][93] = 0;
        pixel_data[105][94] = 0;
        pixel_data[105][95] = 0;
        pixel_data[105][96] = 0;
        pixel_data[105][97] = 0;
        pixel_data[105][98] = 0;
        pixel_data[105][99] = 0;
        pixel_data[105][100] = 0;
        pixel_data[105][101] = 0;
        pixel_data[105][102] = 0;
        pixel_data[105][103] = 0;
        pixel_data[105][104] = 0;
        pixel_data[105][105] = 0;
        pixel_data[105][106] = 0;
        pixel_data[105][107] = 0;
        pixel_data[105][108] = 0;
        pixel_data[105][109] = 0;
        pixel_data[105][110] = 0;
        pixel_data[105][111] = 0;
        pixel_data[105][112] = 0;
        pixel_data[105][113] = 0;
        pixel_data[105][114] = 0;
        pixel_data[105][115] = 0;
        pixel_data[105][116] = 0;
        pixel_data[105][117] = 0;
        pixel_data[105][118] = 0;
        pixel_data[105][119] = 0;
        pixel_data[105][120] = 0;
        pixel_data[105][121] = 0;
        pixel_data[105][122] = 0;
        pixel_data[105][123] = 0;
        pixel_data[105][124] = 0;
        pixel_data[105][125] = 0;
        pixel_data[105][126] = 0;
        pixel_data[105][127] = 0;
        pixel_data[105][128] = 0;
        pixel_data[105][129] = 0;
        pixel_data[105][130] = 0;
        pixel_data[105][131] = 0;
        pixel_data[105][132] = 0;
        pixel_data[105][133] = 0;
        pixel_data[105][134] = 0;
        pixel_data[105][135] = 0;
        pixel_data[105][136] = 0;
        pixel_data[105][137] = 0;
        pixel_data[105][138] = 0;
        pixel_data[105][139] = 0;
        pixel_data[105][140] = 0;
        pixel_data[105][141] = 0;
        pixel_data[105][142] = 0;
        pixel_data[105][143] = 0;
        pixel_data[105][144] = 0;
        pixel_data[105][145] = 0;
        pixel_data[105][146] = 0;
        pixel_data[105][147] = 0;
        pixel_data[105][148] = 0;
        pixel_data[105][149] = 0;
        pixel_data[105][150] = 0;
        pixel_data[105][151] = 0;
        pixel_data[105][152] = 0;
        pixel_data[105][153] = 0;
        pixel_data[105][154] = 0;
        pixel_data[105][155] = 0;
        pixel_data[105][156] = 0;
        pixel_data[105][157] = 0;
        pixel_data[105][158] = 0;
        pixel_data[105][159] = 0;
        pixel_data[105][160] = 0;
        pixel_data[105][161] = 0;
        pixel_data[105][162] = 0;
        pixel_data[105][163] = 0;
        pixel_data[105][164] = 0;
        pixel_data[105][165] = 0;
        pixel_data[105][166] = 0;
        pixel_data[105][167] = 0;
        pixel_data[105][168] = 0;
        pixel_data[105][169] = 0;
        pixel_data[105][170] = 0;
        pixel_data[105][171] = 0;
        pixel_data[105][172] = 0;
        pixel_data[105][173] = 0;
        pixel_data[105][174] = 0;
        pixel_data[105][175] = 0;
        pixel_data[105][176] = 0;
        pixel_data[105][177] = 0;
        pixel_data[105][178] = 0;
        pixel_data[105][179] = 0;
        pixel_data[105][180] = 0;
        pixel_data[105][181] = 0;
        pixel_data[105][182] = 0;
        pixel_data[105][183] = 0;
        pixel_data[105][184] = 0;
        pixel_data[105][185] = 0;
        pixel_data[105][186] = 0;
        pixel_data[105][187] = 0;
        pixel_data[105][188] = 0;
        pixel_data[105][189] = 0;
        pixel_data[105][190] = 0;
        pixel_data[105][191] = 0;
        pixel_data[105][192] = 0;
        pixel_data[105][193] = 0;
        pixel_data[105][194] = 0;
        pixel_data[105][195] = 0;
        pixel_data[105][196] = 0;
        pixel_data[105][197] = 0;
        pixel_data[105][198] = 0;
        pixel_data[105][199] = 0; // y=105
        pixel_data[106][0] = 0;
        pixel_data[106][1] = 0;
        pixel_data[106][2] = 0;
        pixel_data[106][3] = 0;
        pixel_data[106][4] = 0;
        pixel_data[106][5] = 0;
        pixel_data[106][6] = 0;
        pixel_data[106][7] = 0;
        pixel_data[106][8] = 0;
        pixel_data[106][9] = 0;
        pixel_data[106][10] = 0;
        pixel_data[106][11] = 0;
        pixel_data[106][12] = 0;
        pixel_data[106][13] = 0;
        pixel_data[106][14] = 0;
        pixel_data[106][15] = 0;
        pixel_data[106][16] = 0;
        pixel_data[106][17] = 0;
        pixel_data[106][18] = 0;
        pixel_data[106][19] = 0;
        pixel_data[106][20] = 0;
        pixel_data[106][21] = 0;
        pixel_data[106][22] = 0;
        pixel_data[106][23] = 0;
        pixel_data[106][24] = 0;
        pixel_data[106][25] = 0;
        pixel_data[106][26] = 0;
        pixel_data[106][27] = 0;
        pixel_data[106][28] = 0;
        pixel_data[106][29] = 0;
        pixel_data[106][30] = 0;
        pixel_data[106][31] = 0;
        pixel_data[106][32] = 0;
        pixel_data[106][33] = 0;
        pixel_data[106][34] = 0;
        pixel_data[106][35] = 0;
        pixel_data[106][36] = 0;
        pixel_data[106][37] = 0;
        pixel_data[106][38] = 0;
        pixel_data[106][39] = 0;
        pixel_data[106][40] = 0;
        pixel_data[106][41] = 0;
        pixel_data[106][42] = 0;
        pixel_data[106][43] = 0;
        pixel_data[106][44] = 0;
        pixel_data[106][45] = 0;
        pixel_data[106][46] = 0;
        pixel_data[106][47] = 0;
        pixel_data[106][48] = 0;
        pixel_data[106][49] = 0;
        pixel_data[106][50] = 0;
        pixel_data[106][51] = 0;
        pixel_data[106][52] = 0;
        pixel_data[106][53] = 0;
        pixel_data[106][54] = 0;
        pixel_data[106][55] = 0;
        pixel_data[106][56] = 0;
        pixel_data[106][57] = 0;
        pixel_data[106][58] = 0;
        pixel_data[106][59] = 0;
        pixel_data[106][60] = 0;
        pixel_data[106][61] = 0;
        pixel_data[106][62] = 0;
        pixel_data[106][63] = 0;
        pixel_data[106][64] = 0;
        pixel_data[106][65] = 0;
        pixel_data[106][66] = 0;
        pixel_data[106][67] = 0;
        pixel_data[106][68] = 0;
        pixel_data[106][69] = 0;
        pixel_data[106][70] = 0;
        pixel_data[106][71] = 0;
        pixel_data[106][72] = 0;
        pixel_data[106][73] = 0;
        pixel_data[106][74] = 0;
        pixel_data[106][75] = 0;
        pixel_data[106][76] = 0;
        pixel_data[106][77] = 0;
        pixel_data[106][78] = 0;
        pixel_data[106][79] = 0;
        pixel_data[106][80] = 0;
        pixel_data[106][81] = 0;
        pixel_data[106][82] = 0;
        pixel_data[106][83] = 0;
        pixel_data[106][84] = 0;
        pixel_data[106][85] = 0;
        pixel_data[106][86] = 0;
        pixel_data[106][87] = 0;
        pixel_data[106][88] = 0;
        pixel_data[106][89] = 0;
        pixel_data[106][90] = 0;
        pixel_data[106][91] = 0;
        pixel_data[106][92] = 0;
        pixel_data[106][93] = 0;
        pixel_data[106][94] = 0;
        pixel_data[106][95] = 0;
        pixel_data[106][96] = 0;
        pixel_data[106][97] = 0;
        pixel_data[106][98] = 0;
        pixel_data[106][99] = 0;
        pixel_data[106][100] = 0;
        pixel_data[106][101] = 0;
        pixel_data[106][102] = 0;
        pixel_data[106][103] = 0;
        pixel_data[106][104] = 0;
        pixel_data[106][105] = 0;
        pixel_data[106][106] = 0;
        pixel_data[106][107] = 0;
        pixel_data[106][108] = 0;
        pixel_data[106][109] = 0;
        pixel_data[106][110] = 0;
        pixel_data[106][111] = 0;
        pixel_data[106][112] = 0;
        pixel_data[106][113] = 0;
        pixel_data[106][114] = 0;
        pixel_data[106][115] = 0;
        pixel_data[106][116] = 0;
        pixel_data[106][117] = 0;
        pixel_data[106][118] = 0;
        pixel_data[106][119] = 0;
        pixel_data[106][120] = 0;
        pixel_data[106][121] = 0;
        pixel_data[106][122] = 0;
        pixel_data[106][123] = 0;
        pixel_data[106][124] = 0;
        pixel_data[106][125] = 0;
        pixel_data[106][126] = 0;
        pixel_data[106][127] = 0;
        pixel_data[106][128] = 0;
        pixel_data[106][129] = 0;
        pixel_data[106][130] = 0;
        pixel_data[106][131] = 0;
        pixel_data[106][132] = 0;
        pixel_data[106][133] = 0;
        pixel_data[106][134] = 0;
        pixel_data[106][135] = 0;
        pixel_data[106][136] = 0;
        pixel_data[106][137] = 0;
        pixel_data[106][138] = 0;
        pixel_data[106][139] = 0;
        pixel_data[106][140] = 0;
        pixel_data[106][141] = 0;
        pixel_data[106][142] = 0;
        pixel_data[106][143] = 0;
        pixel_data[106][144] = 0;
        pixel_data[106][145] = 0;
        pixel_data[106][146] = 0;
        pixel_data[106][147] = 0;
        pixel_data[106][148] = 0;
        pixel_data[106][149] = 0;
        pixel_data[106][150] = 0;
        pixel_data[106][151] = 0;
        pixel_data[106][152] = 0;
        pixel_data[106][153] = 0;
        pixel_data[106][154] = 0;
        pixel_data[106][155] = 0;
        pixel_data[106][156] = 0;
        pixel_data[106][157] = 0;
        pixel_data[106][158] = 0;
        pixel_data[106][159] = 0;
        pixel_data[106][160] = 0;
        pixel_data[106][161] = 0;
        pixel_data[106][162] = 0;
        pixel_data[106][163] = 0;
        pixel_data[106][164] = 0;
        pixel_data[106][165] = 0;
        pixel_data[106][166] = 0;
        pixel_data[106][167] = 0;
        pixel_data[106][168] = 0;
        pixel_data[106][169] = 0;
        pixel_data[106][170] = 0;
        pixel_data[106][171] = 0;
        pixel_data[106][172] = 0;
        pixel_data[106][173] = 0;
        pixel_data[106][174] = 0;
        pixel_data[106][175] = 0;
        pixel_data[106][176] = 0;
        pixel_data[106][177] = 0;
        pixel_data[106][178] = 0;
        pixel_data[106][179] = 0;
        pixel_data[106][180] = 0;
        pixel_data[106][181] = 0;
        pixel_data[106][182] = 0;
        pixel_data[106][183] = 0;
        pixel_data[106][184] = 0;
        pixel_data[106][185] = 0;
        pixel_data[106][186] = 0;
        pixel_data[106][187] = 0;
        pixel_data[106][188] = 0;
        pixel_data[106][189] = 0;
        pixel_data[106][190] = 0;
        pixel_data[106][191] = 0;
        pixel_data[106][192] = 0;
        pixel_data[106][193] = 0;
        pixel_data[106][194] = 0;
        pixel_data[106][195] = 0;
        pixel_data[106][196] = 0;
        pixel_data[106][197] = 0;
        pixel_data[106][198] = 0;
        pixel_data[106][199] = 0; // y=106
        pixel_data[107][0] = 0;
        pixel_data[107][1] = 0;
        pixel_data[107][2] = 0;
        pixel_data[107][3] = 0;
        pixel_data[107][4] = 0;
        pixel_data[107][5] = 0;
        pixel_data[107][6] = 0;
        pixel_data[107][7] = 0;
        pixel_data[107][8] = 0;
        pixel_data[107][9] = 0;
        pixel_data[107][10] = 0;
        pixel_data[107][11] = 0;
        pixel_data[107][12] = 0;
        pixel_data[107][13] = 0;
        pixel_data[107][14] = 0;
        pixel_data[107][15] = 0;
        pixel_data[107][16] = 0;
        pixel_data[107][17] = 0;
        pixel_data[107][18] = 0;
        pixel_data[107][19] = 0;
        pixel_data[107][20] = 0;
        pixel_data[107][21] = 0;
        pixel_data[107][22] = 0;
        pixel_data[107][23] = 0;
        pixel_data[107][24] = 0;
        pixel_data[107][25] = 0;
        pixel_data[107][26] = 0;
        pixel_data[107][27] = 0;
        pixel_data[107][28] = 0;
        pixel_data[107][29] = 0;
        pixel_data[107][30] = 0;
        pixel_data[107][31] = 0;
        pixel_data[107][32] = 0;
        pixel_data[107][33] = 0;
        pixel_data[107][34] = 0;
        pixel_data[107][35] = 0;
        pixel_data[107][36] = 0;
        pixel_data[107][37] = 0;
        pixel_data[107][38] = 0;
        pixel_data[107][39] = 0;
        pixel_data[107][40] = 0;
        pixel_data[107][41] = 0;
        pixel_data[107][42] = 0;
        pixel_data[107][43] = 0;
        pixel_data[107][44] = 0;
        pixel_data[107][45] = 0;
        pixel_data[107][46] = 0;
        pixel_data[107][47] = 0;
        pixel_data[107][48] = 0;
        pixel_data[107][49] = 0;
        pixel_data[107][50] = 0;
        pixel_data[107][51] = 0;
        pixel_data[107][52] = 0;
        pixel_data[107][53] = 0;
        pixel_data[107][54] = 0;
        pixel_data[107][55] = 0;
        pixel_data[107][56] = 0;
        pixel_data[107][57] = 0;
        pixel_data[107][58] = 0;
        pixel_data[107][59] = 0;
        pixel_data[107][60] = 0;
        pixel_data[107][61] = 0;
        pixel_data[107][62] = 0;
        pixel_data[107][63] = 0;
        pixel_data[107][64] = 0;
        pixel_data[107][65] = 0;
        pixel_data[107][66] = 0;
        pixel_data[107][67] = 0;
        pixel_data[107][68] = 0;
        pixel_data[107][69] = 0;
        pixel_data[107][70] = 0;
        pixel_data[107][71] = 0;
        pixel_data[107][72] = 0;
        pixel_data[107][73] = 0;
        pixel_data[107][74] = 0;
        pixel_data[107][75] = 0;
        pixel_data[107][76] = 0;
        pixel_data[107][77] = 0;
        pixel_data[107][78] = 0;
        pixel_data[107][79] = 0;
        pixel_data[107][80] = 0;
        pixel_data[107][81] = 0;
        pixel_data[107][82] = 0;
        pixel_data[107][83] = 0;
        pixel_data[107][84] = 0;
        pixel_data[107][85] = 0;
        pixel_data[107][86] = 0;
        pixel_data[107][87] = 0;
        pixel_data[107][88] = 0;
        pixel_data[107][89] = 0;
        pixel_data[107][90] = 0;
        pixel_data[107][91] = 0;
        pixel_data[107][92] = 0;
        pixel_data[107][93] = 0;
        pixel_data[107][94] = 0;
        pixel_data[107][95] = 0;
        pixel_data[107][96] = 0;
        pixel_data[107][97] = 0;
        pixel_data[107][98] = 0;
        pixel_data[107][99] = 0;
        pixel_data[107][100] = 0;
        pixel_data[107][101] = 0;
        pixel_data[107][102] = 0;
        pixel_data[107][103] = 0;
        pixel_data[107][104] = 0;
        pixel_data[107][105] = 0;
        pixel_data[107][106] = 0;
        pixel_data[107][107] = 0;
        pixel_data[107][108] = 0;
        pixel_data[107][109] = 0;
        pixel_data[107][110] = 0;
        pixel_data[107][111] = 0;
        pixel_data[107][112] = 0;
        pixel_data[107][113] = 0;
        pixel_data[107][114] = 0;
        pixel_data[107][115] = 0;
        pixel_data[107][116] = 0;
        pixel_data[107][117] = 0;
        pixel_data[107][118] = 0;
        pixel_data[107][119] = 0;
        pixel_data[107][120] = 0;
        pixel_data[107][121] = 0;
        pixel_data[107][122] = 0;
        pixel_data[107][123] = 0;
        pixel_data[107][124] = 0;
        pixel_data[107][125] = 0;
        pixel_data[107][126] = 0;
        pixel_data[107][127] = 0;
        pixel_data[107][128] = 0;
        pixel_data[107][129] = 0;
        pixel_data[107][130] = 0;
        pixel_data[107][131] = 0;
        pixel_data[107][132] = 0;
        pixel_data[107][133] = 0;
        pixel_data[107][134] = 0;
        pixel_data[107][135] = 0;
        pixel_data[107][136] = 0;
        pixel_data[107][137] = 0;
        pixel_data[107][138] = 0;
        pixel_data[107][139] = 0;
        pixel_data[107][140] = 0;
        pixel_data[107][141] = 0;
        pixel_data[107][142] = 0;
        pixel_data[107][143] = 0;
        pixel_data[107][144] = 0;
        pixel_data[107][145] = 0;
        pixel_data[107][146] = 0;
        pixel_data[107][147] = 0;
        pixel_data[107][148] = 0;
        pixel_data[107][149] = 0;
        pixel_data[107][150] = 0;
        pixel_data[107][151] = 0;
        pixel_data[107][152] = 0;
        pixel_data[107][153] = 0;
        pixel_data[107][154] = 0;
        pixel_data[107][155] = 0;
        pixel_data[107][156] = 0;
        pixel_data[107][157] = 0;
        pixel_data[107][158] = 0;
        pixel_data[107][159] = 0;
        pixel_data[107][160] = 0;
        pixel_data[107][161] = 0;
        pixel_data[107][162] = 0;
        pixel_data[107][163] = 0;
        pixel_data[107][164] = 0;
        pixel_data[107][165] = 0;
        pixel_data[107][166] = 0;
        pixel_data[107][167] = 0;
        pixel_data[107][168] = 0;
        pixel_data[107][169] = 0;
        pixel_data[107][170] = 0;
        pixel_data[107][171] = 0;
        pixel_data[107][172] = 0;
        pixel_data[107][173] = 0;
        pixel_data[107][174] = 0;
        pixel_data[107][175] = 0;
        pixel_data[107][176] = 0;
        pixel_data[107][177] = 0;
        pixel_data[107][178] = 0;
        pixel_data[107][179] = 0;
        pixel_data[107][180] = 0;
        pixel_data[107][181] = 0;
        pixel_data[107][182] = 0;
        pixel_data[107][183] = 0;
        pixel_data[107][184] = 0;
        pixel_data[107][185] = 0;
        pixel_data[107][186] = 0;
        pixel_data[107][187] = 0;
        pixel_data[107][188] = 0;
        pixel_data[107][189] = 0;
        pixel_data[107][190] = 0;
        pixel_data[107][191] = 0;
        pixel_data[107][192] = 0;
        pixel_data[107][193] = 0;
        pixel_data[107][194] = 0;
        pixel_data[107][195] = 0;
        pixel_data[107][196] = 0;
        pixel_data[107][197] = 0;
        pixel_data[107][198] = 0;
        pixel_data[107][199] = 0; // y=107
        pixel_data[108][0] = 0;
        pixel_data[108][1] = 0;
        pixel_data[108][2] = 0;
        pixel_data[108][3] = 0;
        pixel_data[108][4] = 0;
        pixel_data[108][5] = 0;
        pixel_data[108][6] = 0;
        pixel_data[108][7] = 0;
        pixel_data[108][8] = 0;
        pixel_data[108][9] = 0;
        pixel_data[108][10] = 0;
        pixel_data[108][11] = 0;
        pixel_data[108][12] = 0;
        pixel_data[108][13] = 0;
        pixel_data[108][14] = 0;
        pixel_data[108][15] = 0;
        pixel_data[108][16] = 0;
        pixel_data[108][17] = 0;
        pixel_data[108][18] = 0;
        pixel_data[108][19] = 0;
        pixel_data[108][20] = 0;
        pixel_data[108][21] = 0;
        pixel_data[108][22] = 0;
        pixel_data[108][23] = 0;
        pixel_data[108][24] = 0;
        pixel_data[108][25] = 0;
        pixel_data[108][26] = 0;
        pixel_data[108][27] = 0;
        pixel_data[108][28] = 0;
        pixel_data[108][29] = 0;
        pixel_data[108][30] = 0;
        pixel_data[108][31] = 0;
        pixel_data[108][32] = 0;
        pixel_data[108][33] = 0;
        pixel_data[108][34] = 0;
        pixel_data[108][35] = 0;
        pixel_data[108][36] = 0;
        pixel_data[108][37] = 0;
        pixel_data[108][38] = 0;
        pixel_data[108][39] = 0;
        pixel_data[108][40] = 0;
        pixel_data[108][41] = 0;
        pixel_data[108][42] = 0;
        pixel_data[108][43] = 0;
        pixel_data[108][44] = 0;
        pixel_data[108][45] = 0;
        pixel_data[108][46] = 0;
        pixel_data[108][47] = 0;
        pixel_data[108][48] = 0;
        pixel_data[108][49] = 0;
        pixel_data[108][50] = 0;
        pixel_data[108][51] = 0;
        pixel_data[108][52] = 0;
        pixel_data[108][53] = 0;
        pixel_data[108][54] = 0;
        pixel_data[108][55] = 0;
        pixel_data[108][56] = 0;
        pixel_data[108][57] = 0;
        pixel_data[108][58] = 0;
        pixel_data[108][59] = 0;
        pixel_data[108][60] = 0;
        pixel_data[108][61] = 0;
        pixel_data[108][62] = 0;
        pixel_data[108][63] = 0;
        pixel_data[108][64] = 0;
        pixel_data[108][65] = 0;
        pixel_data[108][66] = 0;
        pixel_data[108][67] = 0;
        pixel_data[108][68] = 0;
        pixel_data[108][69] = 0;
        pixel_data[108][70] = 0;
        pixel_data[108][71] = 0;
        pixel_data[108][72] = 0;
        pixel_data[108][73] = 0;
        pixel_data[108][74] = 0;
        pixel_data[108][75] = 0;
        pixel_data[108][76] = 0;
        pixel_data[108][77] = 0;
        pixel_data[108][78] = 0;
        pixel_data[108][79] = 0;
        pixel_data[108][80] = 0;
        pixel_data[108][81] = 0;
        pixel_data[108][82] = 0;
        pixel_data[108][83] = 0;
        pixel_data[108][84] = 0;
        pixel_data[108][85] = 0;
        pixel_data[108][86] = 0;
        pixel_data[108][87] = 0;
        pixel_data[108][88] = 0;
        pixel_data[108][89] = 0;
        pixel_data[108][90] = 0;
        pixel_data[108][91] = 0;
        pixel_data[108][92] = 0;
        pixel_data[108][93] = 0;
        pixel_data[108][94] = 0;
        pixel_data[108][95] = 0;
        pixel_data[108][96] = 0;
        pixel_data[108][97] = 0;
        pixel_data[108][98] = 0;
        pixel_data[108][99] = 0;
        pixel_data[108][100] = 0;
        pixel_data[108][101] = 0;
        pixel_data[108][102] = 0;
        pixel_data[108][103] = 0;
        pixel_data[108][104] = 0;
        pixel_data[108][105] = 0;
        pixel_data[108][106] = 0;
        pixel_data[108][107] = 0;
        pixel_data[108][108] = 0;
        pixel_data[108][109] = 0;
        pixel_data[108][110] = 0;
        pixel_data[108][111] = 0;
        pixel_data[108][112] = 0;
        pixel_data[108][113] = 0;
        pixel_data[108][114] = 0;
        pixel_data[108][115] = 0;
        pixel_data[108][116] = 0;
        pixel_data[108][117] = 0;
        pixel_data[108][118] = 0;
        pixel_data[108][119] = 0;
        pixel_data[108][120] = 0;
        pixel_data[108][121] = 0;
        pixel_data[108][122] = 0;
        pixel_data[108][123] = 0;
        pixel_data[108][124] = 0;
        pixel_data[108][125] = 0;
        pixel_data[108][126] = 0;
        pixel_data[108][127] = 0;
        pixel_data[108][128] = 0;
        pixel_data[108][129] = 0;
        pixel_data[108][130] = 0;
        pixel_data[108][131] = 0;
        pixel_data[108][132] = 0;
        pixel_data[108][133] = 0;
        pixel_data[108][134] = 0;
        pixel_data[108][135] = 0;
        pixel_data[108][136] = 0;
        pixel_data[108][137] = 0;
        pixel_data[108][138] = 0;
        pixel_data[108][139] = 0;
        pixel_data[108][140] = 0;
        pixel_data[108][141] = 0;
        pixel_data[108][142] = 0;
        pixel_data[108][143] = 0;
        pixel_data[108][144] = 0;
        pixel_data[108][145] = 0;
        pixel_data[108][146] = 0;
        pixel_data[108][147] = 0;
        pixel_data[108][148] = 0;
        pixel_data[108][149] = 0;
        pixel_data[108][150] = 0;
        pixel_data[108][151] = 0;
        pixel_data[108][152] = 0;
        pixel_data[108][153] = 0;
        pixel_data[108][154] = 0;
        pixel_data[108][155] = 0;
        pixel_data[108][156] = 0;
        pixel_data[108][157] = 0;
        pixel_data[108][158] = 0;
        pixel_data[108][159] = 0;
        pixel_data[108][160] = 0;
        pixel_data[108][161] = 0;
        pixel_data[108][162] = 0;
        pixel_data[108][163] = 0;
        pixel_data[108][164] = 0;
        pixel_data[108][165] = 0;
        pixel_data[108][166] = 0;
        pixel_data[108][167] = 0;
        pixel_data[108][168] = 0;
        pixel_data[108][169] = 0;
        pixel_data[108][170] = 0;
        pixel_data[108][171] = 0;
        pixel_data[108][172] = 0;
        pixel_data[108][173] = 0;
        pixel_data[108][174] = 0;
        pixel_data[108][175] = 0;
        pixel_data[108][176] = 0;
        pixel_data[108][177] = 0;
        pixel_data[108][178] = 0;
        pixel_data[108][179] = 0;
        pixel_data[108][180] = 0;
        pixel_data[108][181] = 0;
        pixel_data[108][182] = 0;
        pixel_data[108][183] = 0;
        pixel_data[108][184] = 0;
        pixel_data[108][185] = 0;
        pixel_data[108][186] = 0;
        pixel_data[108][187] = 0;
        pixel_data[108][188] = 0;
        pixel_data[108][189] = 0;
        pixel_data[108][190] = 0;
        pixel_data[108][191] = 0;
        pixel_data[108][192] = 0;
        pixel_data[108][193] = 0;
        pixel_data[108][194] = 0;
        pixel_data[108][195] = 0;
        pixel_data[108][196] = 0;
        pixel_data[108][197] = 0;
        pixel_data[108][198] = 0;
        pixel_data[108][199] = 0; // y=108
        pixel_data[109][0] = 0;
        pixel_data[109][1] = 0;
        pixel_data[109][2] = 0;
        pixel_data[109][3] = 0;
        pixel_data[109][4] = 0;
        pixel_data[109][5] = 0;
        pixel_data[109][6] = 0;
        pixel_data[109][7] = 0;
        pixel_data[109][8] = 0;
        pixel_data[109][9] = 0;
        pixel_data[109][10] = 0;
        pixel_data[109][11] = 0;
        pixel_data[109][12] = 0;
        pixel_data[109][13] = 0;
        pixel_data[109][14] = 0;
        pixel_data[109][15] = 0;
        pixel_data[109][16] = 0;
        pixel_data[109][17] = 0;
        pixel_data[109][18] = 0;
        pixel_data[109][19] = 0;
        pixel_data[109][20] = 0;
        pixel_data[109][21] = 0;
        pixel_data[109][22] = 0;
        pixel_data[109][23] = 0;
        pixel_data[109][24] = 0;
        pixel_data[109][25] = 0;
        pixel_data[109][26] = 0;
        pixel_data[109][27] = 0;
        pixel_data[109][28] = 0;
        pixel_data[109][29] = 0;
        pixel_data[109][30] = 0;
        pixel_data[109][31] = 0;
        pixel_data[109][32] = 0;
        pixel_data[109][33] = 0;
        pixel_data[109][34] = 0;
        pixel_data[109][35] = 0;
        pixel_data[109][36] = 0;
        pixel_data[109][37] = 0;
        pixel_data[109][38] = 0;
        pixel_data[109][39] = 0;
        pixel_data[109][40] = 0;
        pixel_data[109][41] = 0;
        pixel_data[109][42] = 0;
        pixel_data[109][43] = 0;
        pixel_data[109][44] = 0;
        pixel_data[109][45] = 0;
        pixel_data[109][46] = 0;
        pixel_data[109][47] = 0;
        pixel_data[109][48] = 0;
        pixel_data[109][49] = 0;
        pixel_data[109][50] = 0;
        pixel_data[109][51] = 0;
        pixel_data[109][52] = 0;
        pixel_data[109][53] = 0;
        pixel_data[109][54] = 0;
        pixel_data[109][55] = 0;
        pixel_data[109][56] = 0;
        pixel_data[109][57] = 0;
        pixel_data[109][58] = 0;
        pixel_data[109][59] = 0;
        pixel_data[109][60] = 0;
        pixel_data[109][61] = 0;
        pixel_data[109][62] = 0;
        pixel_data[109][63] = 0;
        pixel_data[109][64] = 0;
        pixel_data[109][65] = 0;
        pixel_data[109][66] = 0;
        pixel_data[109][67] = 0;
        pixel_data[109][68] = 0;
        pixel_data[109][69] = 0;
        pixel_data[109][70] = 0;
        pixel_data[109][71] = 0;
        pixel_data[109][72] = 0;
        pixel_data[109][73] = 0;
        pixel_data[109][74] = 0;
        pixel_data[109][75] = 0;
        pixel_data[109][76] = 0;
        pixel_data[109][77] = 0;
        pixel_data[109][78] = 0;
        pixel_data[109][79] = 0;
        pixel_data[109][80] = 0;
        pixel_data[109][81] = 0;
        pixel_data[109][82] = 0;
        pixel_data[109][83] = 0;
        pixel_data[109][84] = 0;
        pixel_data[109][85] = 0;
        pixel_data[109][86] = 0;
        pixel_data[109][87] = 0;
        pixel_data[109][88] = 0;
        pixel_data[109][89] = 0;
        pixel_data[109][90] = 0;
        pixel_data[109][91] = 0;
        pixel_data[109][92] = 0;
        pixel_data[109][93] = 0;
        pixel_data[109][94] = 0;
        pixel_data[109][95] = 0;
        pixel_data[109][96] = 0;
        pixel_data[109][97] = 0;
        pixel_data[109][98] = 0;
        pixel_data[109][99] = 0;
        pixel_data[109][100] = 0;
        pixel_data[109][101] = 0;
        pixel_data[109][102] = 0;
        pixel_data[109][103] = 0;
        pixel_data[109][104] = 0;
        pixel_data[109][105] = 0;
        pixel_data[109][106] = 0;
        pixel_data[109][107] = 0;
        pixel_data[109][108] = 0;
        pixel_data[109][109] = 0;
        pixel_data[109][110] = 0;
        pixel_data[109][111] = 0;
        pixel_data[109][112] = 0;
        pixel_data[109][113] = 0;
        pixel_data[109][114] = 0;
        pixel_data[109][115] = 0;
        pixel_data[109][116] = 0;
        pixel_data[109][117] = 0;
        pixel_data[109][118] = 0;
        pixel_data[109][119] = 0;
        pixel_data[109][120] = 0;
        pixel_data[109][121] = 0;
        pixel_data[109][122] = 0;
        pixel_data[109][123] = 0;
        pixel_data[109][124] = 0;
        pixel_data[109][125] = 0;
        pixel_data[109][126] = 0;
        pixel_data[109][127] = 0;
        pixel_data[109][128] = 0;
        pixel_data[109][129] = 0;
        pixel_data[109][130] = 0;
        pixel_data[109][131] = 0;
        pixel_data[109][132] = 0;
        pixel_data[109][133] = 0;
        pixel_data[109][134] = 0;
        pixel_data[109][135] = 0;
        pixel_data[109][136] = 0;
        pixel_data[109][137] = 0;
        pixel_data[109][138] = 0;
        pixel_data[109][139] = 0;
        pixel_data[109][140] = 0;
        pixel_data[109][141] = 0;
        pixel_data[109][142] = 0;
        pixel_data[109][143] = 0;
        pixel_data[109][144] = 0;
        pixel_data[109][145] = 0;
        pixel_data[109][146] = 0;
        pixel_data[109][147] = 0;
        pixel_data[109][148] = 0;
        pixel_data[109][149] = 0;
        pixel_data[109][150] = 0;
        pixel_data[109][151] = 0;
        pixel_data[109][152] = 0;
        pixel_data[109][153] = 0;
        pixel_data[109][154] = 0;
        pixel_data[109][155] = 0;
        pixel_data[109][156] = 0;
        pixel_data[109][157] = 0;
        pixel_data[109][158] = 0;
        pixel_data[109][159] = 0;
        pixel_data[109][160] = 0;
        pixel_data[109][161] = 0;
        pixel_data[109][162] = 0;
        pixel_data[109][163] = 0;
        pixel_data[109][164] = 0;
        pixel_data[109][165] = 0;
        pixel_data[109][166] = 0;
        pixel_data[109][167] = 0;
        pixel_data[109][168] = 0;
        pixel_data[109][169] = 0;
        pixel_data[109][170] = 0;
        pixel_data[109][171] = 0;
        pixel_data[109][172] = 0;
        pixel_data[109][173] = 0;
        pixel_data[109][174] = 0;
        pixel_data[109][175] = 0;
        pixel_data[109][176] = 0;
        pixel_data[109][177] = 0;
        pixel_data[109][178] = 0;
        pixel_data[109][179] = 0;
        pixel_data[109][180] = 0;
        pixel_data[109][181] = 0;
        pixel_data[109][182] = 0;
        pixel_data[109][183] = 0;
        pixel_data[109][184] = 0;
        pixel_data[109][185] = 0;
        pixel_data[109][186] = 0;
        pixel_data[109][187] = 0;
        pixel_data[109][188] = 0;
        pixel_data[109][189] = 0;
        pixel_data[109][190] = 0;
        pixel_data[109][191] = 0;
        pixel_data[109][192] = 0;
        pixel_data[109][193] = 0;
        pixel_data[109][194] = 0;
        pixel_data[109][195] = 0;
        pixel_data[109][196] = 0;
        pixel_data[109][197] = 0;
        pixel_data[109][198] = 0;
        pixel_data[109][199] = 0; // y=109
        pixel_data[110][0] = 0;
        pixel_data[110][1] = 0;
        pixel_data[110][2] = 0;
        pixel_data[110][3] = 0;
        pixel_data[110][4] = 0;
        pixel_data[110][5] = 0;
        pixel_data[110][6] = 0;
        pixel_data[110][7] = 0;
        pixel_data[110][8] = 0;
        pixel_data[110][9] = 0;
        pixel_data[110][10] = 0;
        pixel_data[110][11] = 0;
        pixel_data[110][12] = 0;
        pixel_data[110][13] = 0;
        pixel_data[110][14] = 0;
        pixel_data[110][15] = 0;
        pixel_data[110][16] = 0;
        pixel_data[110][17] = 0;
        pixel_data[110][18] = 0;
        pixel_data[110][19] = 0;
        pixel_data[110][20] = 0;
        pixel_data[110][21] = 0;
        pixel_data[110][22] = 0;
        pixel_data[110][23] = 0;
        pixel_data[110][24] = 0;
        pixel_data[110][25] = 0;
        pixel_data[110][26] = 0;
        pixel_data[110][27] = 0;
        pixel_data[110][28] = 0;
        pixel_data[110][29] = 0;
        pixel_data[110][30] = 0;
        pixel_data[110][31] = 0;
        pixel_data[110][32] = 0;
        pixel_data[110][33] = 0;
        pixel_data[110][34] = 0;
        pixel_data[110][35] = 0;
        pixel_data[110][36] = 0;
        pixel_data[110][37] = 0;
        pixel_data[110][38] = 0;
        pixel_data[110][39] = 0;
        pixel_data[110][40] = 0;
        pixel_data[110][41] = 0;
        pixel_data[110][42] = 0;
        pixel_data[110][43] = 0;
        pixel_data[110][44] = 0;
        pixel_data[110][45] = 0;
        pixel_data[110][46] = 0;
        pixel_data[110][47] = 0;
        pixel_data[110][48] = 0;
        pixel_data[110][49] = 0;
        pixel_data[110][50] = 0;
        pixel_data[110][51] = 0;
        pixel_data[110][52] = 0;
        pixel_data[110][53] = 0;
        pixel_data[110][54] = 0;
        pixel_data[110][55] = 0;
        pixel_data[110][56] = 0;
        pixel_data[110][57] = 0;
        pixel_data[110][58] = 0;
        pixel_data[110][59] = 0;
        pixel_data[110][60] = 0;
        pixel_data[110][61] = 0;
        pixel_data[110][62] = 0;
        pixel_data[110][63] = 0;
        pixel_data[110][64] = 0;
        pixel_data[110][65] = 0;
        pixel_data[110][66] = 0;
        pixel_data[110][67] = 0;
        pixel_data[110][68] = 0;
        pixel_data[110][69] = 0;
        pixel_data[110][70] = 0;
        pixel_data[110][71] = 0;
        pixel_data[110][72] = 0;
        pixel_data[110][73] = 0;
        pixel_data[110][74] = 0;
        pixel_data[110][75] = 0;
        pixel_data[110][76] = 0;
        pixel_data[110][77] = 0;
        pixel_data[110][78] = 0;
        pixel_data[110][79] = 0;
        pixel_data[110][80] = 0;
        pixel_data[110][81] = 0;
        pixel_data[110][82] = 0;
        pixel_data[110][83] = 0;
        pixel_data[110][84] = 0;
        pixel_data[110][85] = 0;
        pixel_data[110][86] = 0;
        pixel_data[110][87] = 0;
        pixel_data[110][88] = 0;
        pixel_data[110][89] = 0;
        pixel_data[110][90] = 0;
        pixel_data[110][91] = 0;
        pixel_data[110][92] = 0;
        pixel_data[110][93] = 0;
        pixel_data[110][94] = 0;
        pixel_data[110][95] = 0;
        pixel_data[110][96] = 0;
        pixel_data[110][97] = 0;
        pixel_data[110][98] = 0;
        pixel_data[110][99] = 0;
        pixel_data[110][100] = 0;
        pixel_data[110][101] = 0;
        pixel_data[110][102] = 0;
        pixel_data[110][103] = 0;
        pixel_data[110][104] = 0;
        pixel_data[110][105] = 0;
        pixel_data[110][106] = 0;
        pixel_data[110][107] = 0;
        pixel_data[110][108] = 0;
        pixel_data[110][109] = 0;
        pixel_data[110][110] = 0;
        pixel_data[110][111] = 0;
        pixel_data[110][112] = 0;
        pixel_data[110][113] = 0;
        pixel_data[110][114] = 0;
        pixel_data[110][115] = 0;
        pixel_data[110][116] = 0;
        pixel_data[110][117] = 0;
        pixel_data[110][118] = 0;
        pixel_data[110][119] = 0;
        pixel_data[110][120] = 0;
        pixel_data[110][121] = 0;
        pixel_data[110][122] = 0;
        pixel_data[110][123] = 0;
        pixel_data[110][124] = 0;
        pixel_data[110][125] = 0;
        pixel_data[110][126] = 0;
        pixel_data[110][127] = 0;
        pixel_data[110][128] = 0;
        pixel_data[110][129] = 0;
        pixel_data[110][130] = 0;
        pixel_data[110][131] = 0;
        pixel_data[110][132] = 0;
        pixel_data[110][133] = 0;
        pixel_data[110][134] = 0;
        pixel_data[110][135] = 0;
        pixel_data[110][136] = 0;
        pixel_data[110][137] = 0;
        pixel_data[110][138] = 0;
        pixel_data[110][139] = 0;
        pixel_data[110][140] = 0;
        pixel_data[110][141] = 0;
        pixel_data[110][142] = 0;
        pixel_data[110][143] = 0;
        pixel_data[110][144] = 0;
        pixel_data[110][145] = 0;
        pixel_data[110][146] = 0;
        pixel_data[110][147] = 0;
        pixel_data[110][148] = 0;
        pixel_data[110][149] = 0;
        pixel_data[110][150] = 0;
        pixel_data[110][151] = 0;
        pixel_data[110][152] = 0;
        pixel_data[110][153] = 0;
        pixel_data[110][154] = 0;
        pixel_data[110][155] = 0;
        pixel_data[110][156] = 0;
        pixel_data[110][157] = 0;
        pixel_data[110][158] = 0;
        pixel_data[110][159] = 0;
        pixel_data[110][160] = 0;
        pixel_data[110][161] = 0;
        pixel_data[110][162] = 0;
        pixel_data[110][163] = 0;
        pixel_data[110][164] = 0;
        pixel_data[110][165] = 0;
        pixel_data[110][166] = 0;
        pixel_data[110][167] = 0;
        pixel_data[110][168] = 0;
        pixel_data[110][169] = 0;
        pixel_data[110][170] = 0;
        pixel_data[110][171] = 0;
        pixel_data[110][172] = 0;
        pixel_data[110][173] = 0;
        pixel_data[110][174] = 0;
        pixel_data[110][175] = 0;
        pixel_data[110][176] = 0;
        pixel_data[110][177] = 0;
        pixel_data[110][178] = 0;
        pixel_data[110][179] = 0;
        pixel_data[110][180] = 0;
        pixel_data[110][181] = 0;
        pixel_data[110][182] = 0;
        pixel_data[110][183] = 0;
        pixel_data[110][184] = 0;
        pixel_data[110][185] = 0;
        pixel_data[110][186] = 0;
        pixel_data[110][187] = 0;
        pixel_data[110][188] = 0;
        pixel_data[110][189] = 0;
        pixel_data[110][190] = 0;
        pixel_data[110][191] = 0;
        pixel_data[110][192] = 0;
        pixel_data[110][193] = 0;
        pixel_data[110][194] = 0;
        pixel_data[110][195] = 0;
        pixel_data[110][196] = 0;
        pixel_data[110][197] = 0;
        pixel_data[110][198] = 0;
        pixel_data[110][199] = 0; // y=110
        pixel_data[111][0] = 0;
        pixel_data[111][1] = 0;
        pixel_data[111][2] = 0;
        pixel_data[111][3] = 0;
        pixel_data[111][4] = 0;
        pixel_data[111][5] = 0;
        pixel_data[111][6] = 0;
        pixel_data[111][7] = 0;
        pixel_data[111][8] = 0;
        pixel_data[111][9] = 0;
        pixel_data[111][10] = 0;
        pixel_data[111][11] = 0;
        pixel_data[111][12] = 0;
        pixel_data[111][13] = 0;
        pixel_data[111][14] = 0;
        pixel_data[111][15] = 0;
        pixel_data[111][16] = 0;
        pixel_data[111][17] = 0;
        pixel_data[111][18] = 0;
        pixel_data[111][19] = 0;
        pixel_data[111][20] = 0;
        pixel_data[111][21] = 0;
        pixel_data[111][22] = 0;
        pixel_data[111][23] = 0;
        pixel_data[111][24] = 0;
        pixel_data[111][25] = 0;
        pixel_data[111][26] = 0;
        pixel_data[111][27] = 0;
        pixel_data[111][28] = 0;
        pixel_data[111][29] = 0;
        pixel_data[111][30] = 0;
        pixel_data[111][31] = 0;
        pixel_data[111][32] = 0;
        pixel_data[111][33] = 0;
        pixel_data[111][34] = 0;
        pixel_data[111][35] = 0;
        pixel_data[111][36] = 0;
        pixel_data[111][37] = 0;
        pixel_data[111][38] = 0;
        pixel_data[111][39] = 0;
        pixel_data[111][40] = 0;
        pixel_data[111][41] = 0;
        pixel_data[111][42] = 0;
        pixel_data[111][43] = 0;
        pixel_data[111][44] = 0;
        pixel_data[111][45] = 0;
        pixel_data[111][46] = 0;
        pixel_data[111][47] = 0;
        pixel_data[111][48] = 0;
        pixel_data[111][49] = 0;
        pixel_data[111][50] = 0;
        pixel_data[111][51] = 0;
        pixel_data[111][52] = 0;
        pixel_data[111][53] = 0;
        pixel_data[111][54] = 0;
        pixel_data[111][55] = 0;
        pixel_data[111][56] = 0;
        pixel_data[111][57] = 0;
        pixel_data[111][58] = 0;
        pixel_data[111][59] = 0;
        pixel_data[111][60] = 0;
        pixel_data[111][61] = 0;
        pixel_data[111][62] = 0;
        pixel_data[111][63] = 0;
        pixel_data[111][64] = 0;
        pixel_data[111][65] = 0;
        pixel_data[111][66] = 0;
        pixel_data[111][67] = 0;
        pixel_data[111][68] = 0;
        pixel_data[111][69] = 0;
        pixel_data[111][70] = 0;
        pixel_data[111][71] = 0;
        pixel_data[111][72] = 0;
        pixel_data[111][73] = 0;
        pixel_data[111][74] = 0;
        pixel_data[111][75] = 0;
        pixel_data[111][76] = 0;
        pixel_data[111][77] = 0;
        pixel_data[111][78] = 0;
        pixel_data[111][79] = 0;
        pixel_data[111][80] = 0;
        pixel_data[111][81] = 0;
        pixel_data[111][82] = 0;
        pixel_data[111][83] = 0;
        pixel_data[111][84] = 0;
        pixel_data[111][85] = 0;
        pixel_data[111][86] = 0;
        pixel_data[111][87] = 0;
        pixel_data[111][88] = 0;
        pixel_data[111][89] = 0;
        pixel_data[111][90] = 0;
        pixel_data[111][91] = 0;
        pixel_data[111][92] = 0;
        pixel_data[111][93] = 0;
        pixel_data[111][94] = 0;
        pixel_data[111][95] = 0;
        pixel_data[111][96] = 0;
        pixel_data[111][97] = 0;
        pixel_data[111][98] = 0;
        pixel_data[111][99] = 0;
        pixel_data[111][100] = 0;
        pixel_data[111][101] = 0;
        pixel_data[111][102] = 0;
        pixel_data[111][103] = 0;
        pixel_data[111][104] = 0;
        pixel_data[111][105] = 0;
        pixel_data[111][106] = 0;
        pixel_data[111][107] = 0;
        pixel_data[111][108] = 0;
        pixel_data[111][109] = 0;
        pixel_data[111][110] = 0;
        pixel_data[111][111] = 0;
        pixel_data[111][112] = 0;
        pixel_data[111][113] = 0;
        pixel_data[111][114] = 0;
        pixel_data[111][115] = 0;
        pixel_data[111][116] = 0;
        pixel_data[111][117] = 0;
        pixel_data[111][118] = 0;
        pixel_data[111][119] = 0;
        pixel_data[111][120] = 0;
        pixel_data[111][121] = 0;
        pixel_data[111][122] = 0;
        pixel_data[111][123] = 0;
        pixel_data[111][124] = 0;
        pixel_data[111][125] = 0;
        pixel_data[111][126] = 0;
        pixel_data[111][127] = 0;
        pixel_data[111][128] = 0;
        pixel_data[111][129] = 0;
        pixel_data[111][130] = 0;
        pixel_data[111][131] = 0;
        pixel_data[111][132] = 0;
        pixel_data[111][133] = 0;
        pixel_data[111][134] = 0;
        pixel_data[111][135] = 0;
        pixel_data[111][136] = 0;
        pixel_data[111][137] = 0;
        pixel_data[111][138] = 0;
        pixel_data[111][139] = 0;
        pixel_data[111][140] = 0;
        pixel_data[111][141] = 0;
        pixel_data[111][142] = 0;
        pixel_data[111][143] = 0;
        pixel_data[111][144] = 0;
        pixel_data[111][145] = 0;
        pixel_data[111][146] = 0;
        pixel_data[111][147] = 0;
        pixel_data[111][148] = 0;
        pixel_data[111][149] = 0;
        pixel_data[111][150] = 0;
        pixel_data[111][151] = 0;
        pixel_data[111][152] = 0;
        pixel_data[111][153] = 0;
        pixel_data[111][154] = 0;
        pixel_data[111][155] = 0;
        pixel_data[111][156] = 0;
        pixel_data[111][157] = 0;
        pixel_data[111][158] = 0;
        pixel_data[111][159] = 0;
        pixel_data[111][160] = 0;
        pixel_data[111][161] = 0;
        pixel_data[111][162] = 0;
        pixel_data[111][163] = 0;
        pixel_data[111][164] = 0;
        pixel_data[111][165] = 0;
        pixel_data[111][166] = 0;
        pixel_data[111][167] = 0;
        pixel_data[111][168] = 0;
        pixel_data[111][169] = 0;
        pixel_data[111][170] = 0;
        pixel_data[111][171] = 0;
        pixel_data[111][172] = 0;
        pixel_data[111][173] = 0;
        pixel_data[111][174] = 0;
        pixel_data[111][175] = 0;
        pixel_data[111][176] = 0;
        pixel_data[111][177] = 0;
        pixel_data[111][178] = 0;
        pixel_data[111][179] = 0;
        pixel_data[111][180] = 0;
        pixel_data[111][181] = 0;
        pixel_data[111][182] = 0;
        pixel_data[111][183] = 0;
        pixel_data[111][184] = 0;
        pixel_data[111][185] = 0;
        pixel_data[111][186] = 0;
        pixel_data[111][187] = 0;
        pixel_data[111][188] = 0;
        pixel_data[111][189] = 0;
        pixel_data[111][190] = 0;
        pixel_data[111][191] = 0;
        pixel_data[111][192] = 0;
        pixel_data[111][193] = 0;
        pixel_data[111][194] = 0;
        pixel_data[111][195] = 0;
        pixel_data[111][196] = 0;
        pixel_data[111][197] = 0;
        pixel_data[111][198] = 0;
        pixel_data[111][199] = 0; // y=111
        pixel_data[112][0] = 0;
        pixel_data[112][1] = 0;
        pixel_data[112][2] = 0;
        pixel_data[112][3] = 0;
        pixel_data[112][4] = 0;
        pixel_data[112][5] = 0;
        pixel_data[112][6] = 0;
        pixel_data[112][7] = 0;
        pixel_data[112][8] = 0;
        pixel_data[112][9] = 0;
        pixel_data[112][10] = 0;
        pixel_data[112][11] = 0;
        pixel_data[112][12] = 0;
        pixel_data[112][13] = 0;
        pixel_data[112][14] = 0;
        pixel_data[112][15] = 0;
        pixel_data[112][16] = 0;
        pixel_data[112][17] = 0;
        pixel_data[112][18] = 0;
        pixel_data[112][19] = 0;
        pixel_data[112][20] = 0;
        pixel_data[112][21] = 0;
        pixel_data[112][22] = 0;
        pixel_data[112][23] = 0;
        pixel_data[112][24] = 0;
        pixel_data[112][25] = 0;
        pixel_data[112][26] = 0;
        pixel_data[112][27] = 0;
        pixel_data[112][28] = 0;
        pixel_data[112][29] = 0;
        pixel_data[112][30] = 0;
        pixel_data[112][31] = 0;
        pixel_data[112][32] = 0;
        pixel_data[112][33] = 0;
        pixel_data[112][34] = 0;
        pixel_data[112][35] = 0;
        pixel_data[112][36] = 0;
        pixel_data[112][37] = 0;
        pixel_data[112][38] = 0;
        pixel_data[112][39] = 0;
        pixel_data[112][40] = 0;
        pixel_data[112][41] = 0;
        pixel_data[112][42] = 0;
        pixel_data[112][43] = 0;
        pixel_data[112][44] = 0;
        pixel_data[112][45] = 0;
        pixel_data[112][46] = 0;
        pixel_data[112][47] = 0;
        pixel_data[112][48] = 0;
        pixel_data[112][49] = 0;
        pixel_data[112][50] = 0;
        pixel_data[112][51] = 0;
        pixel_data[112][52] = 0;
        pixel_data[112][53] = 0;
        pixel_data[112][54] = 0;
        pixel_data[112][55] = 0;
        pixel_data[112][56] = 0;
        pixel_data[112][57] = 0;
        pixel_data[112][58] = 0;
        pixel_data[112][59] = 0;
        pixel_data[112][60] = 0;
        pixel_data[112][61] = 0;
        pixel_data[112][62] = 0;
        pixel_data[112][63] = 0;
        pixel_data[112][64] = 0;
        pixel_data[112][65] = 0;
        pixel_data[112][66] = 0;
        pixel_data[112][67] = 0;
        pixel_data[112][68] = 0;
        pixel_data[112][69] = 0;
        pixel_data[112][70] = 0;
        pixel_data[112][71] = 0;
        pixel_data[112][72] = 0;
        pixel_data[112][73] = 0;
        pixel_data[112][74] = 0;
        pixel_data[112][75] = 0;
        pixel_data[112][76] = 0;
        pixel_data[112][77] = 0;
        pixel_data[112][78] = 0;
        pixel_data[112][79] = 0;
        pixel_data[112][80] = 0;
        pixel_data[112][81] = 0;
        pixel_data[112][82] = 0;
        pixel_data[112][83] = 0;
        pixel_data[112][84] = 0;
        pixel_data[112][85] = 0;
        pixel_data[112][86] = 0;
        pixel_data[112][87] = 0;
        pixel_data[112][88] = 0;
        pixel_data[112][89] = 0;
        pixel_data[112][90] = 0;
        pixel_data[112][91] = 0;
        pixel_data[112][92] = 0;
        pixel_data[112][93] = 0;
        pixel_data[112][94] = 0;
        pixel_data[112][95] = 0;
        pixel_data[112][96] = 0;
        pixel_data[112][97] = 0;
        pixel_data[112][98] = 0;
        pixel_data[112][99] = 0;
        pixel_data[112][100] = 0;
        pixel_data[112][101] = 0;
        pixel_data[112][102] = 0;
        pixel_data[112][103] = 0;
        pixel_data[112][104] = 0;
        pixel_data[112][105] = 0;
        pixel_data[112][106] = 0;
        pixel_data[112][107] = 0;
        pixel_data[112][108] = 0;
        pixel_data[112][109] = 0;
        pixel_data[112][110] = 0;
        pixel_data[112][111] = 0;
        pixel_data[112][112] = 0;
        pixel_data[112][113] = 0;
        pixel_data[112][114] = 0;
        pixel_data[112][115] = 0;
        pixel_data[112][116] = 0;
        pixel_data[112][117] = 0;
        pixel_data[112][118] = 0;
        pixel_data[112][119] = 0;
        pixel_data[112][120] = 0;
        pixel_data[112][121] = 0;
        pixel_data[112][122] = 0;
        pixel_data[112][123] = 0;
        pixel_data[112][124] = 0;
        pixel_data[112][125] = 0;
        pixel_data[112][126] = 0;
        pixel_data[112][127] = 0;
        pixel_data[112][128] = 0;
        pixel_data[112][129] = 0;
        pixel_data[112][130] = 0;
        pixel_data[112][131] = 0;
        pixel_data[112][132] = 0;
        pixel_data[112][133] = 0;
        pixel_data[112][134] = 0;
        pixel_data[112][135] = 0;
        pixel_data[112][136] = 0;
        pixel_data[112][137] = 0;
        pixel_data[112][138] = 0;
        pixel_data[112][139] = 0;
        pixel_data[112][140] = 0;
        pixel_data[112][141] = 0;
        pixel_data[112][142] = 0;
        pixel_data[112][143] = 0;
        pixel_data[112][144] = 0;
        pixel_data[112][145] = 0;
        pixel_data[112][146] = 0;
        pixel_data[112][147] = 0;
        pixel_data[112][148] = 0;
        pixel_data[112][149] = 0;
        pixel_data[112][150] = 0;
        pixel_data[112][151] = 0;
        pixel_data[112][152] = 0;
        pixel_data[112][153] = 0;
        pixel_data[112][154] = 0;
        pixel_data[112][155] = 0;
        pixel_data[112][156] = 0;
        pixel_data[112][157] = 0;
        pixel_data[112][158] = 0;
        pixel_data[112][159] = 0;
        pixel_data[112][160] = 0;
        pixel_data[112][161] = 0;
        pixel_data[112][162] = 0;
        pixel_data[112][163] = 0;
        pixel_data[112][164] = 0;
        pixel_data[112][165] = 0;
        pixel_data[112][166] = 0;
        pixel_data[112][167] = 0;
        pixel_data[112][168] = 0;
        pixel_data[112][169] = 0;
        pixel_data[112][170] = 0;
        pixel_data[112][171] = 0;
        pixel_data[112][172] = 0;
        pixel_data[112][173] = 0;
        pixel_data[112][174] = 0;
        pixel_data[112][175] = 0;
        pixel_data[112][176] = 0;
        pixel_data[112][177] = 0;
        pixel_data[112][178] = 0;
        pixel_data[112][179] = 0;
        pixel_data[112][180] = 0;
        pixel_data[112][181] = 0;
        pixel_data[112][182] = 0;
        pixel_data[112][183] = 0;
        pixel_data[112][184] = 0;
        pixel_data[112][185] = 0;
        pixel_data[112][186] = 0;
        pixel_data[112][187] = 0;
        pixel_data[112][188] = 0;
        pixel_data[112][189] = 0;
        pixel_data[112][190] = 0;
        pixel_data[112][191] = 0;
        pixel_data[112][192] = 0;
        pixel_data[112][193] = 0;
        pixel_data[112][194] = 0;
        pixel_data[112][195] = 0;
        pixel_data[112][196] = 0;
        pixel_data[112][197] = 0;
        pixel_data[112][198] = 0;
        pixel_data[112][199] = 0; // y=112
        pixel_data[113][0] = 0;
        pixel_data[113][1] = 0;
        pixel_data[113][2] = 0;
        pixel_data[113][3] = 0;
        pixel_data[113][4] = 0;
        pixel_data[113][5] = 0;
        pixel_data[113][6] = 0;
        pixel_data[113][7] = 0;
        pixel_data[113][8] = 0;
        pixel_data[113][9] = 0;
        pixel_data[113][10] = 0;
        pixel_data[113][11] = 0;
        pixel_data[113][12] = 0;
        pixel_data[113][13] = 0;
        pixel_data[113][14] = 0;
        pixel_data[113][15] = 0;
        pixel_data[113][16] = 0;
        pixel_data[113][17] = 0;
        pixel_data[113][18] = 0;
        pixel_data[113][19] = 0;
        pixel_data[113][20] = 0;
        pixel_data[113][21] = 0;
        pixel_data[113][22] = 0;
        pixel_data[113][23] = 0;
        pixel_data[113][24] = 0;
        pixel_data[113][25] = 0;
        pixel_data[113][26] = 0;
        pixel_data[113][27] = 0;
        pixel_data[113][28] = 0;
        pixel_data[113][29] = 0;
        pixel_data[113][30] = 0;
        pixel_data[113][31] = 0;
        pixel_data[113][32] = 0;
        pixel_data[113][33] = 0;
        pixel_data[113][34] = 0;
        pixel_data[113][35] = 0;
        pixel_data[113][36] = 0;
        pixel_data[113][37] = 0;
        pixel_data[113][38] = 0;
        pixel_data[113][39] = 0;
        pixel_data[113][40] = 0;
        pixel_data[113][41] = 0;
        pixel_data[113][42] = 0;
        pixel_data[113][43] = 0;
        pixel_data[113][44] = 0;
        pixel_data[113][45] = 0;
        pixel_data[113][46] = 0;
        pixel_data[113][47] = 0;
        pixel_data[113][48] = 0;
        pixel_data[113][49] = 0;
        pixel_data[113][50] = 0;
        pixel_data[113][51] = 0;
        pixel_data[113][52] = 0;
        pixel_data[113][53] = 0;
        pixel_data[113][54] = 0;
        pixel_data[113][55] = 0;
        pixel_data[113][56] = 0;
        pixel_data[113][57] = 0;
        pixel_data[113][58] = 0;
        pixel_data[113][59] = 0;
        pixel_data[113][60] = 0;
        pixel_data[113][61] = 0;
        pixel_data[113][62] = 0;
        pixel_data[113][63] = 0;
        pixel_data[113][64] = 0;
        pixel_data[113][65] = 0;
        pixel_data[113][66] = 0;
        pixel_data[113][67] = 0;
        pixel_data[113][68] = 0;
        pixel_data[113][69] = 0;
        pixel_data[113][70] = 0;
        pixel_data[113][71] = 0;
        pixel_data[113][72] = 0;
        pixel_data[113][73] = 0;
        pixel_data[113][74] = 0;
        pixel_data[113][75] = 0;
        pixel_data[113][76] = 0;
        pixel_data[113][77] = 0;
        pixel_data[113][78] = 0;
        pixel_data[113][79] = 0;
        pixel_data[113][80] = 0;
        pixel_data[113][81] = 0;
        pixel_data[113][82] = 0;
        pixel_data[113][83] = 0;
        pixel_data[113][84] = 0;
        pixel_data[113][85] = 0;
        pixel_data[113][86] = 0;
        pixel_data[113][87] = 0;
        pixel_data[113][88] = 0;
        pixel_data[113][89] = 0;
        pixel_data[113][90] = 0;
        pixel_data[113][91] = 0;
        pixel_data[113][92] = 0;
        pixel_data[113][93] = 0;
        pixel_data[113][94] = 0;
        pixel_data[113][95] = 0;
        pixel_data[113][96] = 0;
        pixel_data[113][97] = 0;
        pixel_data[113][98] = 0;
        pixel_data[113][99] = 0;
        pixel_data[113][100] = 0;
        pixel_data[113][101] = 0;
        pixel_data[113][102] = 0;
        pixel_data[113][103] = 0;
        pixel_data[113][104] = 0;
        pixel_data[113][105] = 0;
        pixel_data[113][106] = 0;
        pixel_data[113][107] = 0;
        pixel_data[113][108] = 0;
        pixel_data[113][109] = 0;
        pixel_data[113][110] = 0;
        pixel_data[113][111] = 0;
        pixel_data[113][112] = 0;
        pixel_data[113][113] = 0;
        pixel_data[113][114] = 0;
        pixel_data[113][115] = 0;
        pixel_data[113][116] = 0;
        pixel_data[113][117] = 0;
        pixel_data[113][118] = 0;
        pixel_data[113][119] = 0;
        pixel_data[113][120] = 0;
        pixel_data[113][121] = 0;
        pixel_data[113][122] = 0;
        pixel_data[113][123] = 0;
        pixel_data[113][124] = 0;
        pixel_data[113][125] = 0;
        pixel_data[113][126] = 0;
        pixel_data[113][127] = 0;
        pixel_data[113][128] = 0;
        pixel_data[113][129] = 0;
        pixel_data[113][130] = 0;
        pixel_data[113][131] = 0;
        pixel_data[113][132] = 0;
        pixel_data[113][133] = 0;
        pixel_data[113][134] = 0;
        pixel_data[113][135] = 0;
        pixel_data[113][136] = 0;
        pixel_data[113][137] = 0;
        pixel_data[113][138] = 0;
        pixel_data[113][139] = 0;
        pixel_data[113][140] = 0;
        pixel_data[113][141] = 0;
        pixel_data[113][142] = 0;
        pixel_data[113][143] = 0;
        pixel_data[113][144] = 0;
        pixel_data[113][145] = 0;
        pixel_data[113][146] = 0;
        pixel_data[113][147] = 0;
        pixel_data[113][148] = 0;
        pixel_data[113][149] = 0;
        pixel_data[113][150] = 0;
        pixel_data[113][151] = 0;
        pixel_data[113][152] = 0;
        pixel_data[113][153] = 0;
        pixel_data[113][154] = 0;
        pixel_data[113][155] = 0;
        pixel_data[113][156] = 0;
        pixel_data[113][157] = 0;
        pixel_data[113][158] = 0;
        pixel_data[113][159] = 0;
        pixel_data[113][160] = 0;
        pixel_data[113][161] = 0;
        pixel_data[113][162] = 0;
        pixel_data[113][163] = 0;
        pixel_data[113][164] = 0;
        pixel_data[113][165] = 0;
        pixel_data[113][166] = 0;
        pixel_data[113][167] = 0;
        pixel_data[113][168] = 0;
        pixel_data[113][169] = 0;
        pixel_data[113][170] = 0;
        pixel_data[113][171] = 0;
        pixel_data[113][172] = 0;
        pixel_data[113][173] = 0;
        pixel_data[113][174] = 0;
        pixel_data[113][175] = 0;
        pixel_data[113][176] = 0;
        pixel_data[113][177] = 0;
        pixel_data[113][178] = 0;
        pixel_data[113][179] = 0;
        pixel_data[113][180] = 0;
        pixel_data[113][181] = 0;
        pixel_data[113][182] = 0;
        pixel_data[113][183] = 0;
        pixel_data[113][184] = 0;
        pixel_data[113][185] = 0;
        pixel_data[113][186] = 0;
        pixel_data[113][187] = 0;
        pixel_data[113][188] = 0;
        pixel_data[113][189] = 0;
        pixel_data[113][190] = 0;
        pixel_data[113][191] = 0;
        pixel_data[113][192] = 0;
        pixel_data[113][193] = 0;
        pixel_data[113][194] = 0;
        pixel_data[113][195] = 0;
        pixel_data[113][196] = 0;
        pixel_data[113][197] = 0;
        pixel_data[113][198] = 0;
        pixel_data[113][199] = 0; // y=113
        pixel_data[114][0] = 0;
        pixel_data[114][1] = 0;
        pixel_data[114][2] = 0;
        pixel_data[114][3] = 0;
        pixel_data[114][4] = 0;
        pixel_data[114][5] = 0;
        pixel_data[114][6] = 0;
        pixel_data[114][7] = 0;
        pixel_data[114][8] = 0;
        pixel_data[114][9] = 0;
        pixel_data[114][10] = 0;
        pixel_data[114][11] = 0;
        pixel_data[114][12] = 0;
        pixel_data[114][13] = 0;
        pixel_data[114][14] = 0;
        pixel_data[114][15] = 0;
        pixel_data[114][16] = 0;
        pixel_data[114][17] = 0;
        pixel_data[114][18] = 0;
        pixel_data[114][19] = 0;
        pixel_data[114][20] = 0;
        pixel_data[114][21] = 0;
        pixel_data[114][22] = 0;
        pixel_data[114][23] = 0;
        pixel_data[114][24] = 0;
        pixel_data[114][25] = 0;
        pixel_data[114][26] = 0;
        pixel_data[114][27] = 0;
        pixel_data[114][28] = 0;
        pixel_data[114][29] = 0;
        pixel_data[114][30] = 0;
        pixel_data[114][31] = 0;
        pixel_data[114][32] = 0;
        pixel_data[114][33] = 0;
        pixel_data[114][34] = 0;
        pixel_data[114][35] = 0;
        pixel_data[114][36] = 0;
        pixel_data[114][37] = 0;
        pixel_data[114][38] = 0;
        pixel_data[114][39] = 0;
        pixel_data[114][40] = 0;
        pixel_data[114][41] = 0;
        pixel_data[114][42] = 0;
        pixel_data[114][43] = 0;
        pixel_data[114][44] = 0;
        pixel_data[114][45] = 0;
        pixel_data[114][46] = 0;
        pixel_data[114][47] = 0;
        pixel_data[114][48] = 0;
        pixel_data[114][49] = 0;
        pixel_data[114][50] = 0;
        pixel_data[114][51] = 0;
        pixel_data[114][52] = 0;
        pixel_data[114][53] = 0;
        pixel_data[114][54] = 0;
        pixel_data[114][55] = 0;
        pixel_data[114][56] = 0;
        pixel_data[114][57] = 0;
        pixel_data[114][58] = 0;
        pixel_data[114][59] = 0;
        pixel_data[114][60] = 0;
        pixel_data[114][61] = 0;
        pixel_data[114][62] = 0;
        pixel_data[114][63] = 0;
        pixel_data[114][64] = 0;
        pixel_data[114][65] = 0;
        pixel_data[114][66] = 0;
        pixel_data[114][67] = 0;
        pixel_data[114][68] = 0;
        pixel_data[114][69] = 0;
        pixel_data[114][70] = 0;
        pixel_data[114][71] = 0;
        pixel_data[114][72] = 0;
        pixel_data[114][73] = 0;
        pixel_data[114][74] = 0;
        pixel_data[114][75] = 0;
        pixel_data[114][76] = 0;
        pixel_data[114][77] = 0;
        pixel_data[114][78] = 0;
        pixel_data[114][79] = 0;
        pixel_data[114][80] = 0;
        pixel_data[114][81] = 0;
        pixel_data[114][82] = 0;
        pixel_data[114][83] = 0;
        pixel_data[114][84] = 0;
        pixel_data[114][85] = 0;
        pixel_data[114][86] = 0;
        pixel_data[114][87] = 0;
        pixel_data[114][88] = 0;
        pixel_data[114][89] = 0;
        pixel_data[114][90] = 0;
        pixel_data[114][91] = 0;
        pixel_data[114][92] = 0;
        pixel_data[114][93] = 0;
        pixel_data[114][94] = 0;
        pixel_data[114][95] = 0;
        pixel_data[114][96] = 0;
        pixel_data[114][97] = 0;
        pixel_data[114][98] = 0;
        pixel_data[114][99] = 0;
        pixel_data[114][100] = 0;
        pixel_data[114][101] = 0;
        pixel_data[114][102] = 0;
        pixel_data[114][103] = 0;
        pixel_data[114][104] = 0;
        pixel_data[114][105] = 0;
        pixel_data[114][106] = 0;
        pixel_data[114][107] = 0;
        pixel_data[114][108] = 0;
        pixel_data[114][109] = 0;
        pixel_data[114][110] = 0;
        pixel_data[114][111] = 0;
        pixel_data[114][112] = 0;
        pixel_data[114][113] = 0;
        pixel_data[114][114] = 0;
        pixel_data[114][115] = 0;
        pixel_data[114][116] = 0;
        pixel_data[114][117] = 0;
        pixel_data[114][118] = 0;
        pixel_data[114][119] = 0;
        pixel_data[114][120] = 0;
        pixel_data[114][121] = 0;
        pixel_data[114][122] = 0;
        pixel_data[114][123] = 0;
        pixel_data[114][124] = 0;
        pixel_data[114][125] = 0;
        pixel_data[114][126] = 0;
        pixel_data[114][127] = 0;
        pixel_data[114][128] = 0;
        pixel_data[114][129] = 0;
        pixel_data[114][130] = 0;
        pixel_data[114][131] = 0;
        pixel_data[114][132] = 0;
        pixel_data[114][133] = 0;
        pixel_data[114][134] = 0;
        pixel_data[114][135] = 0;
        pixel_data[114][136] = 0;
        pixel_data[114][137] = 0;
        pixel_data[114][138] = 0;
        pixel_data[114][139] = 0;
        pixel_data[114][140] = 0;
        pixel_data[114][141] = 0;
        pixel_data[114][142] = 0;
        pixel_data[114][143] = 0;
        pixel_data[114][144] = 0;
        pixel_data[114][145] = 0;
        pixel_data[114][146] = 0;
        pixel_data[114][147] = 0;
        pixel_data[114][148] = 0;
        pixel_data[114][149] = 0;
        pixel_data[114][150] = 0;
        pixel_data[114][151] = 0;
        pixel_data[114][152] = 0;
        pixel_data[114][153] = 0;
        pixel_data[114][154] = 0;
        pixel_data[114][155] = 0;
        pixel_data[114][156] = 0;
        pixel_data[114][157] = 0;
        pixel_data[114][158] = 0;
        pixel_data[114][159] = 0;
        pixel_data[114][160] = 0;
        pixel_data[114][161] = 0;
        pixel_data[114][162] = 0;
        pixel_data[114][163] = 0;
        pixel_data[114][164] = 0;
        pixel_data[114][165] = 0;
        pixel_data[114][166] = 0;
        pixel_data[114][167] = 0;
        pixel_data[114][168] = 0;
        pixel_data[114][169] = 0;
        pixel_data[114][170] = 0;
        pixel_data[114][171] = 0;
        pixel_data[114][172] = 0;
        pixel_data[114][173] = 0;
        pixel_data[114][174] = 0;
        pixel_data[114][175] = 0;
        pixel_data[114][176] = 0;
        pixel_data[114][177] = 0;
        pixel_data[114][178] = 0;
        pixel_data[114][179] = 0;
        pixel_data[114][180] = 0;
        pixel_data[114][181] = 0;
        pixel_data[114][182] = 0;
        pixel_data[114][183] = 0;
        pixel_data[114][184] = 0;
        pixel_data[114][185] = 0;
        pixel_data[114][186] = 0;
        pixel_data[114][187] = 0;
        pixel_data[114][188] = 0;
        pixel_data[114][189] = 0;
        pixel_data[114][190] = 0;
        pixel_data[114][191] = 0;
        pixel_data[114][192] = 0;
        pixel_data[114][193] = 0;
        pixel_data[114][194] = 0;
        pixel_data[114][195] = 0;
        pixel_data[114][196] = 0;
        pixel_data[114][197] = 0;
        pixel_data[114][198] = 0;
        pixel_data[114][199] = 0; // y=114
        pixel_data[115][0] = 0;
        pixel_data[115][1] = 0;
        pixel_data[115][2] = 0;
        pixel_data[115][3] = 0;
        pixel_data[115][4] = 0;
        pixel_data[115][5] = 0;
        pixel_data[115][6] = 0;
        pixel_data[115][7] = 0;
        pixel_data[115][8] = 0;
        pixel_data[115][9] = 0;
        pixel_data[115][10] = 0;
        pixel_data[115][11] = 0;
        pixel_data[115][12] = 0;
        pixel_data[115][13] = 0;
        pixel_data[115][14] = 0;
        pixel_data[115][15] = 0;
        pixel_data[115][16] = 0;
        pixel_data[115][17] = 0;
        pixel_data[115][18] = 0;
        pixel_data[115][19] = 0;
        pixel_data[115][20] = 0;
        pixel_data[115][21] = 0;
        pixel_data[115][22] = 0;
        pixel_data[115][23] = 0;
        pixel_data[115][24] = 0;
        pixel_data[115][25] = 0;
        pixel_data[115][26] = 0;
        pixel_data[115][27] = 0;
        pixel_data[115][28] = 0;
        pixel_data[115][29] = 0;
        pixel_data[115][30] = 0;
        pixel_data[115][31] = 0;
        pixel_data[115][32] = 0;
        pixel_data[115][33] = 0;
        pixel_data[115][34] = 0;
        pixel_data[115][35] = 0;
        pixel_data[115][36] = 0;
        pixel_data[115][37] = 0;
        pixel_data[115][38] = 0;
        pixel_data[115][39] = 0;
        pixel_data[115][40] = 0;
        pixel_data[115][41] = 0;
        pixel_data[115][42] = 0;
        pixel_data[115][43] = 0;
        pixel_data[115][44] = 0;
        pixel_data[115][45] = 0;
        pixel_data[115][46] = 0;
        pixel_data[115][47] = 0;
        pixel_data[115][48] = 0;
        pixel_data[115][49] = 0;
        pixel_data[115][50] = 0;
        pixel_data[115][51] = 0;
        pixel_data[115][52] = 0;
        pixel_data[115][53] = 0;
        pixel_data[115][54] = 0;
        pixel_data[115][55] = 0;
        pixel_data[115][56] = 0;
        pixel_data[115][57] = 0;
        pixel_data[115][58] = 0;
        pixel_data[115][59] = 0;
        pixel_data[115][60] = 0;
        pixel_data[115][61] = 0;
        pixel_data[115][62] = 0;
        pixel_data[115][63] = 0;
        pixel_data[115][64] = 0;
        pixel_data[115][65] = 0;
        pixel_data[115][66] = 0;
        pixel_data[115][67] = 0;
        pixel_data[115][68] = 0;
        pixel_data[115][69] = 0;
        pixel_data[115][70] = 0;
        pixel_data[115][71] = 0;
        pixel_data[115][72] = 0;
        pixel_data[115][73] = 0;
        pixel_data[115][74] = 0;
        pixel_data[115][75] = 0;
        pixel_data[115][76] = 0;
        pixel_data[115][77] = 0;
        pixel_data[115][78] = 0;
        pixel_data[115][79] = 0;
        pixel_data[115][80] = 0;
        pixel_data[115][81] = 0;
        pixel_data[115][82] = 0;
        pixel_data[115][83] = 0;
        pixel_data[115][84] = 0;
        pixel_data[115][85] = 0;
        pixel_data[115][86] = 0;
        pixel_data[115][87] = 0;
        pixel_data[115][88] = 0;
        pixel_data[115][89] = 0;
        pixel_data[115][90] = 0;
        pixel_data[115][91] = 0;
        pixel_data[115][92] = 0;
        pixel_data[115][93] = 0;
        pixel_data[115][94] = 0;
        pixel_data[115][95] = 0;
        pixel_data[115][96] = 0;
        pixel_data[115][97] = 0;
        pixel_data[115][98] = 0;
        pixel_data[115][99] = 0;
        pixel_data[115][100] = 0;
        pixel_data[115][101] = 0;
        pixel_data[115][102] = 0;
        pixel_data[115][103] = 0;
        pixel_data[115][104] = 0;
        pixel_data[115][105] = 0;
        pixel_data[115][106] = 0;
        pixel_data[115][107] = 0;
        pixel_data[115][108] = 0;
        pixel_data[115][109] = 0;
        pixel_data[115][110] = 0;
        pixel_data[115][111] = 0;
        pixel_data[115][112] = 0;
        pixel_data[115][113] = 0;
        pixel_data[115][114] = 0;
        pixel_data[115][115] = 0;
        pixel_data[115][116] = 0;
        pixel_data[115][117] = 0;
        pixel_data[115][118] = 0;
        pixel_data[115][119] = 0;
        pixel_data[115][120] = 0;
        pixel_data[115][121] = 0;
        pixel_data[115][122] = 0;
        pixel_data[115][123] = 0;
        pixel_data[115][124] = 0;
        pixel_data[115][125] = 0;
        pixel_data[115][126] = 0;
        pixel_data[115][127] = 0;
        pixel_data[115][128] = 0;
        pixel_data[115][129] = 0;
        pixel_data[115][130] = 0;
        pixel_data[115][131] = 0;
        pixel_data[115][132] = 0;
        pixel_data[115][133] = 0;
        pixel_data[115][134] = 0;
        pixel_data[115][135] = 0;
        pixel_data[115][136] = 0;
        pixel_data[115][137] = 0;
        pixel_data[115][138] = 0;
        pixel_data[115][139] = 0;
        pixel_data[115][140] = 0;
        pixel_data[115][141] = 0;
        pixel_data[115][142] = 0;
        pixel_data[115][143] = 0;
        pixel_data[115][144] = 0;
        pixel_data[115][145] = 0;
        pixel_data[115][146] = 0;
        pixel_data[115][147] = 0;
        pixel_data[115][148] = 0;
        pixel_data[115][149] = 0;
        pixel_data[115][150] = 0;
        pixel_data[115][151] = 0;
        pixel_data[115][152] = 0;
        pixel_data[115][153] = 0;
        pixel_data[115][154] = 0;
        pixel_data[115][155] = 0;
        pixel_data[115][156] = 0;
        pixel_data[115][157] = 0;
        pixel_data[115][158] = 0;
        pixel_data[115][159] = 0;
        pixel_data[115][160] = 0;
        pixel_data[115][161] = 0;
        pixel_data[115][162] = 0;
        pixel_data[115][163] = 0;
        pixel_data[115][164] = 0;
        pixel_data[115][165] = 0;
        pixel_data[115][166] = 0;
        pixel_data[115][167] = 0;
        pixel_data[115][168] = 0;
        pixel_data[115][169] = 0;
        pixel_data[115][170] = 0;
        pixel_data[115][171] = 0;
        pixel_data[115][172] = 0;
        pixel_data[115][173] = 0;
        pixel_data[115][174] = 0;
        pixel_data[115][175] = 0;
        pixel_data[115][176] = 0;
        pixel_data[115][177] = 0;
        pixel_data[115][178] = 0;
        pixel_data[115][179] = 0;
        pixel_data[115][180] = 0;
        pixel_data[115][181] = 0;
        pixel_data[115][182] = 0;
        pixel_data[115][183] = 0;
        pixel_data[115][184] = 0;
        pixel_data[115][185] = 0;
        pixel_data[115][186] = 0;
        pixel_data[115][187] = 0;
        pixel_data[115][188] = 0;
        pixel_data[115][189] = 0;
        pixel_data[115][190] = 0;
        pixel_data[115][191] = 0;
        pixel_data[115][192] = 0;
        pixel_data[115][193] = 0;
        pixel_data[115][194] = 0;
        pixel_data[115][195] = 0;
        pixel_data[115][196] = 0;
        pixel_data[115][197] = 0;
        pixel_data[115][198] = 0;
        pixel_data[115][199] = 0; // y=115
        pixel_data[116][0] = 0;
        pixel_data[116][1] = 0;
        pixel_data[116][2] = 0;
        pixel_data[116][3] = 0;
        pixel_data[116][4] = 0;
        pixel_data[116][5] = 0;
        pixel_data[116][6] = 0;
        pixel_data[116][7] = 0;
        pixel_data[116][8] = 0;
        pixel_data[116][9] = 0;
        pixel_data[116][10] = 0;
        pixel_data[116][11] = 0;
        pixel_data[116][12] = 0;
        pixel_data[116][13] = 0;
        pixel_data[116][14] = 0;
        pixel_data[116][15] = 0;
        pixel_data[116][16] = 0;
        pixel_data[116][17] = 0;
        pixel_data[116][18] = 0;
        pixel_data[116][19] = 0;
        pixel_data[116][20] = 0;
        pixel_data[116][21] = 0;
        pixel_data[116][22] = 0;
        pixel_data[116][23] = 0;
        pixel_data[116][24] = 0;
        pixel_data[116][25] = 0;
        pixel_data[116][26] = 0;
        pixel_data[116][27] = 0;
        pixel_data[116][28] = 0;
        pixel_data[116][29] = 0;
        pixel_data[116][30] = 0;
        pixel_data[116][31] = 0;
        pixel_data[116][32] = 0;
        pixel_data[116][33] = 0;
        pixel_data[116][34] = 0;
        pixel_data[116][35] = 0;
        pixel_data[116][36] = 0;
        pixel_data[116][37] = 0;
        pixel_data[116][38] = 0;
        pixel_data[116][39] = 0;
        pixel_data[116][40] = 0;
        pixel_data[116][41] = 0;
        pixel_data[116][42] = 0;
        pixel_data[116][43] = 0;
        pixel_data[116][44] = 0;
        pixel_data[116][45] = 0;
        pixel_data[116][46] = 0;
        pixel_data[116][47] = 0;
        pixel_data[116][48] = 0;
        pixel_data[116][49] = 0;
        pixel_data[116][50] = 0;
        pixel_data[116][51] = 0;
        pixel_data[116][52] = 0;
        pixel_data[116][53] = 0;
        pixel_data[116][54] = 0;
        pixel_data[116][55] = 0;
        pixel_data[116][56] = 0;
        pixel_data[116][57] = 0;
        pixel_data[116][58] = 0;
        pixel_data[116][59] = 0;
        pixel_data[116][60] = 0;
        pixel_data[116][61] = 0;
        pixel_data[116][62] = 0;
        pixel_data[116][63] = 0;
        pixel_data[116][64] = 0;
        pixel_data[116][65] = 0;
        pixel_data[116][66] = 0;
        pixel_data[116][67] = 0;
        pixel_data[116][68] = 0;
        pixel_data[116][69] = 0;
        pixel_data[116][70] = 0;
        pixel_data[116][71] = 0;
        pixel_data[116][72] = 0;
        pixel_data[116][73] = 0;
        pixel_data[116][74] = 0;
        pixel_data[116][75] = 0;
        pixel_data[116][76] = 0;
        pixel_data[116][77] = 0;
        pixel_data[116][78] = 0;
        pixel_data[116][79] = 0;
        pixel_data[116][80] = 0;
        pixel_data[116][81] = 0;
        pixel_data[116][82] = 0;
        pixel_data[116][83] = 0;
        pixel_data[116][84] = 0;
        pixel_data[116][85] = 0;
        pixel_data[116][86] = 0;
        pixel_data[116][87] = 0;
        pixel_data[116][88] = 0;
        pixel_data[116][89] = 0;
        pixel_data[116][90] = 0;
        pixel_data[116][91] = 0;
        pixel_data[116][92] = 0;
        pixel_data[116][93] = 0;
        pixel_data[116][94] = 0;
        pixel_data[116][95] = 0;
        pixel_data[116][96] = 0;
        pixel_data[116][97] = 0;
        pixel_data[116][98] = 0;
        pixel_data[116][99] = 0;
        pixel_data[116][100] = 0;
        pixel_data[116][101] = 0;
        pixel_data[116][102] = 0;
        pixel_data[116][103] = 0;
        pixel_data[116][104] = 0;
        pixel_data[116][105] = 0;
        pixel_data[116][106] = 0;
        pixel_data[116][107] = 0;
        pixel_data[116][108] = 0;
        pixel_data[116][109] = 0;
        pixel_data[116][110] = 0;
        pixel_data[116][111] = 0;
        pixel_data[116][112] = 0;
        pixel_data[116][113] = 0;
        pixel_data[116][114] = 0;
        pixel_data[116][115] = 0;
        pixel_data[116][116] = 0;
        pixel_data[116][117] = 0;
        pixel_data[116][118] = 0;
        pixel_data[116][119] = 0;
        pixel_data[116][120] = 0;
        pixel_data[116][121] = 0;
        pixel_data[116][122] = 0;
        pixel_data[116][123] = 0;
        pixel_data[116][124] = 0;
        pixel_data[116][125] = 0;
        pixel_data[116][126] = 0;
        pixel_data[116][127] = 0;
        pixel_data[116][128] = 0;
        pixel_data[116][129] = 0;
        pixel_data[116][130] = 0;
        pixel_data[116][131] = 0;
        pixel_data[116][132] = 0;
        pixel_data[116][133] = 0;
        pixel_data[116][134] = 0;
        pixel_data[116][135] = 0;
        pixel_data[116][136] = 0;
        pixel_data[116][137] = 0;
        pixel_data[116][138] = 0;
        pixel_data[116][139] = 0;
        pixel_data[116][140] = 0;
        pixel_data[116][141] = 0;
        pixel_data[116][142] = 0;
        pixel_data[116][143] = 0;
        pixel_data[116][144] = 0;
        pixel_data[116][145] = 0;
        pixel_data[116][146] = 0;
        pixel_data[116][147] = 0;
        pixel_data[116][148] = 0;
        pixel_data[116][149] = 0;
        pixel_data[116][150] = 0;
        pixel_data[116][151] = 0;
        pixel_data[116][152] = 0;
        pixel_data[116][153] = 0;
        pixel_data[116][154] = 0;
        pixel_data[116][155] = 0;
        pixel_data[116][156] = 0;
        pixel_data[116][157] = 0;
        pixel_data[116][158] = 0;
        pixel_data[116][159] = 0;
        pixel_data[116][160] = 0;
        pixel_data[116][161] = 0;
        pixel_data[116][162] = 0;
        pixel_data[116][163] = 0;
        pixel_data[116][164] = 0;
        pixel_data[116][165] = 0;
        pixel_data[116][166] = 0;
        pixel_data[116][167] = 0;
        pixel_data[116][168] = 0;
        pixel_data[116][169] = 0;
        pixel_data[116][170] = 0;
        pixel_data[116][171] = 0;
        pixel_data[116][172] = 0;
        pixel_data[116][173] = 0;
        pixel_data[116][174] = 0;
        pixel_data[116][175] = 0;
        pixel_data[116][176] = 0;
        pixel_data[116][177] = 0;
        pixel_data[116][178] = 0;
        pixel_data[116][179] = 0;
        pixel_data[116][180] = 0;
        pixel_data[116][181] = 0;
        pixel_data[116][182] = 0;
        pixel_data[116][183] = 0;
        pixel_data[116][184] = 0;
        pixel_data[116][185] = 0;
        pixel_data[116][186] = 0;
        pixel_data[116][187] = 0;
        pixel_data[116][188] = 0;
        pixel_data[116][189] = 0;
        pixel_data[116][190] = 0;
        pixel_data[116][191] = 0;
        pixel_data[116][192] = 0;
        pixel_data[116][193] = 0;
        pixel_data[116][194] = 0;
        pixel_data[116][195] = 0;
        pixel_data[116][196] = 0;
        pixel_data[116][197] = 0;
        pixel_data[116][198] = 0;
        pixel_data[116][199] = 0; // y=116
        pixel_data[117][0] = 0;
        pixel_data[117][1] = 0;
        pixel_data[117][2] = 0;
        pixel_data[117][3] = 0;
        pixel_data[117][4] = 0;
        pixel_data[117][5] = 0;
        pixel_data[117][6] = 0;
        pixel_data[117][7] = 0;
        pixel_data[117][8] = 0;
        pixel_data[117][9] = 0;
        pixel_data[117][10] = 0;
        pixel_data[117][11] = 0;
        pixel_data[117][12] = 0;
        pixel_data[117][13] = 0;
        pixel_data[117][14] = 0;
        pixel_data[117][15] = 0;
        pixel_data[117][16] = 0;
        pixel_data[117][17] = 0;
        pixel_data[117][18] = 0;
        pixel_data[117][19] = 0;
        pixel_data[117][20] = 0;
        pixel_data[117][21] = 0;
        pixel_data[117][22] = 0;
        pixel_data[117][23] = 0;
        pixel_data[117][24] = 0;
        pixel_data[117][25] = 0;
        pixel_data[117][26] = 0;
        pixel_data[117][27] = 0;
        pixel_data[117][28] = 0;
        pixel_data[117][29] = 0;
        pixel_data[117][30] = 0;
        pixel_data[117][31] = 0;
        pixel_data[117][32] = 0;
        pixel_data[117][33] = 0;
        pixel_data[117][34] = 0;
        pixel_data[117][35] = 0;
        pixel_data[117][36] = 0;
        pixel_data[117][37] = 0;
        pixel_data[117][38] = 0;
        pixel_data[117][39] = 0;
        pixel_data[117][40] = 0;
        pixel_data[117][41] = 0;
        pixel_data[117][42] = 0;
        pixel_data[117][43] = 0;
        pixel_data[117][44] = 0;
        pixel_data[117][45] = 0;
        pixel_data[117][46] = 0;
        pixel_data[117][47] = 0;
        pixel_data[117][48] = 0;
        pixel_data[117][49] = 0;
        pixel_data[117][50] = 0;
        pixel_data[117][51] = 0;
        pixel_data[117][52] = 0;
        pixel_data[117][53] = 0;
        pixel_data[117][54] = 0;
        pixel_data[117][55] = 0;
        pixel_data[117][56] = 0;
        pixel_data[117][57] = 0;
        pixel_data[117][58] = 0;
        pixel_data[117][59] = 0;
        pixel_data[117][60] = 0;
        pixel_data[117][61] = 0;
        pixel_data[117][62] = 0;
        pixel_data[117][63] = 0;
        pixel_data[117][64] = 0;
        pixel_data[117][65] = 0;
        pixel_data[117][66] = 0;
        pixel_data[117][67] = 0;
        pixel_data[117][68] = 0;
        pixel_data[117][69] = 0;
        pixel_data[117][70] = 0;
        pixel_data[117][71] = 0;
        pixel_data[117][72] = 0;
        pixel_data[117][73] = 0;
        pixel_data[117][74] = 0;
        pixel_data[117][75] = 0;
        pixel_data[117][76] = 0;
        pixel_data[117][77] = 0;
        pixel_data[117][78] = 0;
        pixel_data[117][79] = 0;
        pixel_data[117][80] = 0;
        pixel_data[117][81] = 0;
        pixel_data[117][82] = 0;
        pixel_data[117][83] = 0;
        pixel_data[117][84] = 0;
        pixel_data[117][85] = 0;
        pixel_data[117][86] = 0;
        pixel_data[117][87] = 0;
        pixel_data[117][88] = 0;
        pixel_data[117][89] = 0;
        pixel_data[117][90] = 0;
        pixel_data[117][91] = 0;
        pixel_data[117][92] = 0;
        pixel_data[117][93] = 0;
        pixel_data[117][94] = 0;
        pixel_data[117][95] = 0;
        pixel_data[117][96] = 0;
        pixel_data[117][97] = 0;
        pixel_data[117][98] = 0;
        pixel_data[117][99] = 0;
        pixel_data[117][100] = 0;
        pixel_data[117][101] = 0;
        pixel_data[117][102] = 0;
        pixel_data[117][103] = 0;
        pixel_data[117][104] = 0;
        pixel_data[117][105] = 0;
        pixel_data[117][106] = 0;
        pixel_data[117][107] = 0;
        pixel_data[117][108] = 0;
        pixel_data[117][109] = 0;
        pixel_data[117][110] = 0;
        pixel_data[117][111] = 0;
        pixel_data[117][112] = 0;
        pixel_data[117][113] = 0;
        pixel_data[117][114] = 0;
        pixel_data[117][115] = 0;
        pixel_data[117][116] = 0;
        pixel_data[117][117] = 0;
        pixel_data[117][118] = 0;
        pixel_data[117][119] = 0;
        pixel_data[117][120] = 0;
        pixel_data[117][121] = 0;
        pixel_data[117][122] = 0;
        pixel_data[117][123] = 0;
        pixel_data[117][124] = 0;
        pixel_data[117][125] = 0;
        pixel_data[117][126] = 0;
        pixel_data[117][127] = 0;
        pixel_data[117][128] = 0;
        pixel_data[117][129] = 0;
        pixel_data[117][130] = 0;
        pixel_data[117][131] = 0;
        pixel_data[117][132] = 0;
        pixel_data[117][133] = 0;
        pixel_data[117][134] = 0;
        pixel_data[117][135] = 0;
        pixel_data[117][136] = 0;
        pixel_data[117][137] = 0;
        pixel_data[117][138] = 0;
        pixel_data[117][139] = 0;
        pixel_data[117][140] = 0;
        pixel_data[117][141] = 0;
        pixel_data[117][142] = 0;
        pixel_data[117][143] = 0;
        pixel_data[117][144] = 0;
        pixel_data[117][145] = 0;
        pixel_data[117][146] = 0;
        pixel_data[117][147] = 0;
        pixel_data[117][148] = 0;
        pixel_data[117][149] = 0;
        pixel_data[117][150] = 0;
        pixel_data[117][151] = 0;
        pixel_data[117][152] = 0;
        pixel_data[117][153] = 0;
        pixel_data[117][154] = 0;
        pixel_data[117][155] = 0;
        pixel_data[117][156] = 0;
        pixel_data[117][157] = 0;
        pixel_data[117][158] = 0;
        pixel_data[117][159] = 0;
        pixel_data[117][160] = 0;
        pixel_data[117][161] = 0;
        pixel_data[117][162] = 0;
        pixel_data[117][163] = 0;
        pixel_data[117][164] = 0;
        pixel_data[117][165] = 0;
        pixel_data[117][166] = 0;
        pixel_data[117][167] = 0;
        pixel_data[117][168] = 0;
        pixel_data[117][169] = 0;
        pixel_data[117][170] = 0;
        pixel_data[117][171] = 0;
        pixel_data[117][172] = 0;
        pixel_data[117][173] = 0;
        pixel_data[117][174] = 0;
        pixel_data[117][175] = 0;
        pixel_data[117][176] = 0;
        pixel_data[117][177] = 0;
        pixel_data[117][178] = 0;
        pixel_data[117][179] = 0;
        pixel_data[117][180] = 0;
        pixel_data[117][181] = 0;
        pixel_data[117][182] = 0;
        pixel_data[117][183] = 0;
        pixel_data[117][184] = 0;
        pixel_data[117][185] = 0;
        pixel_data[117][186] = 0;
        pixel_data[117][187] = 0;
        pixel_data[117][188] = 0;
        pixel_data[117][189] = 0;
        pixel_data[117][190] = 0;
        pixel_data[117][191] = 0;
        pixel_data[117][192] = 0;
        pixel_data[117][193] = 0;
        pixel_data[117][194] = 0;
        pixel_data[117][195] = 0;
        pixel_data[117][196] = 0;
        pixel_data[117][197] = 0;
        pixel_data[117][198] = 0;
        pixel_data[117][199] = 0; // y=117
        pixel_data[118][0] = 0;
        pixel_data[118][1] = 0;
        pixel_data[118][2] = 0;
        pixel_data[118][3] = 0;
        pixel_data[118][4] = 0;
        pixel_data[118][5] = 0;
        pixel_data[118][6] = 0;
        pixel_data[118][7] = 0;
        pixel_data[118][8] = 0;
        pixel_data[118][9] = 0;
        pixel_data[118][10] = 0;
        pixel_data[118][11] = 0;
        pixel_data[118][12] = 0;
        pixel_data[118][13] = 0;
        pixel_data[118][14] = 0;
        pixel_data[118][15] = 0;
        pixel_data[118][16] = 0;
        pixel_data[118][17] = 0;
        pixel_data[118][18] = 0;
        pixel_data[118][19] = 0;
        pixel_data[118][20] = 0;
        pixel_data[118][21] = 0;
        pixel_data[118][22] = 0;
        pixel_data[118][23] = 0;
        pixel_data[118][24] = 0;
        pixel_data[118][25] = 0;
        pixel_data[118][26] = 0;
        pixel_data[118][27] = 0;
        pixel_data[118][28] = 0;
        pixel_data[118][29] = 0;
        pixel_data[118][30] = 0;
        pixel_data[118][31] = 0;
        pixel_data[118][32] = 0;
        pixel_data[118][33] = 0;
        pixel_data[118][34] = 0;
        pixel_data[118][35] = 0;
        pixel_data[118][36] = 0;
        pixel_data[118][37] = 0;
        pixel_data[118][38] = 0;
        pixel_data[118][39] = 0;
        pixel_data[118][40] = 0;
        pixel_data[118][41] = 0;
        pixel_data[118][42] = 0;
        pixel_data[118][43] = 0;
        pixel_data[118][44] = 0;
        pixel_data[118][45] = 0;
        pixel_data[118][46] = 0;
        pixel_data[118][47] = 0;
        pixel_data[118][48] = 0;
        pixel_data[118][49] = 0;
        pixel_data[118][50] = 0;
        pixel_data[118][51] = 0;
        pixel_data[118][52] = 0;
        pixel_data[118][53] = 0;
        pixel_data[118][54] = 0;
        pixel_data[118][55] = 0;
        pixel_data[118][56] = 0;
        pixel_data[118][57] = 0;
        pixel_data[118][58] = 0;
        pixel_data[118][59] = 0;
        pixel_data[118][60] = 0;
        pixel_data[118][61] = 0;
        pixel_data[118][62] = 0;
        pixel_data[118][63] = 0;
        pixel_data[118][64] = 0;
        pixel_data[118][65] = 0;
        pixel_data[118][66] = 0;
        pixel_data[118][67] = 0;
        pixel_data[118][68] = 0;
        pixel_data[118][69] = 0;
        pixel_data[118][70] = 0;
        pixel_data[118][71] = 0;
        pixel_data[118][72] = 0;
        pixel_data[118][73] = 0;
        pixel_data[118][74] = 0;
        pixel_data[118][75] = 0;
        pixel_data[118][76] = 0;
        pixel_data[118][77] = 0;
        pixel_data[118][78] = 0;
        pixel_data[118][79] = 0;
        pixel_data[118][80] = 0;
        pixel_data[118][81] = 0;
        pixel_data[118][82] = 0;
        pixel_data[118][83] = 0;
        pixel_data[118][84] = 0;
        pixel_data[118][85] = 0;
        pixel_data[118][86] = 0;
        pixel_data[118][87] = 0;
        pixel_data[118][88] = 0;
        pixel_data[118][89] = 0;
        pixel_data[118][90] = 0;
        pixel_data[118][91] = 0;
        pixel_data[118][92] = 0;
        pixel_data[118][93] = 0;
        pixel_data[118][94] = 0;
        pixel_data[118][95] = 0;
        pixel_data[118][96] = 0;
        pixel_data[118][97] = 0;
        pixel_data[118][98] = 0;
        pixel_data[118][99] = 0;
        pixel_data[118][100] = 0;
        pixel_data[118][101] = 0;
        pixel_data[118][102] = 0;
        pixel_data[118][103] = 0;
        pixel_data[118][104] = 0;
        pixel_data[118][105] = 0;
        pixel_data[118][106] = 0;
        pixel_data[118][107] = 0;
        pixel_data[118][108] = 0;
        pixel_data[118][109] = 0;
        pixel_data[118][110] = 0;
        pixel_data[118][111] = 0;
        pixel_data[118][112] = 0;
        pixel_data[118][113] = 0;
        pixel_data[118][114] = 0;
        pixel_data[118][115] = 0;
        pixel_data[118][116] = 0;
        pixel_data[118][117] = 0;
        pixel_data[118][118] = 0;
        pixel_data[118][119] = 0;
        pixel_data[118][120] = 0;
        pixel_data[118][121] = 0;
        pixel_data[118][122] = 0;
        pixel_data[118][123] = 0;
        pixel_data[118][124] = 0;
        pixel_data[118][125] = 0;
        pixel_data[118][126] = 0;
        pixel_data[118][127] = 0;
        pixel_data[118][128] = 0;
        pixel_data[118][129] = 0;
        pixel_data[118][130] = 0;
        pixel_data[118][131] = 0;
        pixel_data[118][132] = 0;
        pixel_data[118][133] = 0;
        pixel_data[118][134] = 0;
        pixel_data[118][135] = 0;
        pixel_data[118][136] = 0;
        pixel_data[118][137] = 0;
        pixel_data[118][138] = 0;
        pixel_data[118][139] = 0;
        pixel_data[118][140] = 0;
        pixel_data[118][141] = 0;
        pixel_data[118][142] = 0;
        pixel_data[118][143] = 0;
        pixel_data[118][144] = 0;
        pixel_data[118][145] = 0;
        pixel_data[118][146] = 0;
        pixel_data[118][147] = 0;
        pixel_data[118][148] = 0;
        pixel_data[118][149] = 0;
        pixel_data[118][150] = 0;
        pixel_data[118][151] = 0;
        pixel_data[118][152] = 0;
        pixel_data[118][153] = 0;
        pixel_data[118][154] = 0;
        pixel_data[118][155] = 0;
        pixel_data[118][156] = 0;
        pixel_data[118][157] = 0;
        pixel_data[118][158] = 0;
        pixel_data[118][159] = 0;
        pixel_data[118][160] = 0;
        pixel_data[118][161] = 0;
        pixel_data[118][162] = 0;
        pixel_data[118][163] = 0;
        pixel_data[118][164] = 0;
        pixel_data[118][165] = 0;
        pixel_data[118][166] = 0;
        pixel_data[118][167] = 0;
        pixel_data[118][168] = 0;
        pixel_data[118][169] = 0;
        pixel_data[118][170] = 0;
        pixel_data[118][171] = 0;
        pixel_data[118][172] = 0;
        pixel_data[118][173] = 0;
        pixel_data[118][174] = 0;
        pixel_data[118][175] = 0;
        pixel_data[118][176] = 0;
        pixel_data[118][177] = 0;
        pixel_data[118][178] = 0;
        pixel_data[118][179] = 0;
        pixel_data[118][180] = 0;
        pixel_data[118][181] = 0;
        pixel_data[118][182] = 0;
        pixel_data[118][183] = 0;
        pixel_data[118][184] = 0;
        pixel_data[118][185] = 0;
        pixel_data[118][186] = 0;
        pixel_data[118][187] = 0;
        pixel_data[118][188] = 0;
        pixel_data[118][189] = 0;
        pixel_data[118][190] = 0;
        pixel_data[118][191] = 0;
        pixel_data[118][192] = 0;
        pixel_data[118][193] = 0;
        pixel_data[118][194] = 0;
        pixel_data[118][195] = 0;
        pixel_data[118][196] = 0;
        pixel_data[118][197] = 0;
        pixel_data[118][198] = 0;
        pixel_data[118][199] = 0; // y=118
        pixel_data[119][0] = 0;
        pixel_data[119][1] = 0;
        pixel_data[119][2] = 0;
        pixel_data[119][3] = 0;
        pixel_data[119][4] = 0;
        pixel_data[119][5] = 0;
        pixel_data[119][6] = 0;
        pixel_data[119][7] = 0;
        pixel_data[119][8] = 0;
        pixel_data[119][9] = 0;
        pixel_data[119][10] = 0;
        pixel_data[119][11] = 0;
        pixel_data[119][12] = 0;
        pixel_data[119][13] = 0;
        pixel_data[119][14] = 0;
        pixel_data[119][15] = 0;
        pixel_data[119][16] = 0;
        pixel_data[119][17] = 0;
        pixel_data[119][18] = 0;
        pixel_data[119][19] = 0;
        pixel_data[119][20] = 0;
        pixel_data[119][21] = 0;
        pixel_data[119][22] = 0;
        pixel_data[119][23] = 0;
        pixel_data[119][24] = 0;
        pixel_data[119][25] = 0;
        pixel_data[119][26] = 0;
        pixel_data[119][27] = 0;
        pixel_data[119][28] = 0;
        pixel_data[119][29] = 0;
        pixel_data[119][30] = 0;
        pixel_data[119][31] = 0;
        pixel_data[119][32] = 0;
        pixel_data[119][33] = 0;
        pixel_data[119][34] = 0;
        pixel_data[119][35] = 0;
        pixel_data[119][36] = 0;
        pixel_data[119][37] = 0;
        pixel_data[119][38] = 0;
        pixel_data[119][39] = 0;
        pixel_data[119][40] = 0;
        pixel_data[119][41] = 0;
        pixel_data[119][42] = 0;
        pixel_data[119][43] = 0;
        pixel_data[119][44] = 0;
        pixel_data[119][45] = 0;
        pixel_data[119][46] = 0;
        pixel_data[119][47] = 0;
        pixel_data[119][48] = 0;
        pixel_data[119][49] = 0;
        pixel_data[119][50] = 0;
        pixel_data[119][51] = 0;
        pixel_data[119][52] = 0;
        pixel_data[119][53] = 0;
        pixel_data[119][54] = 0;
        pixel_data[119][55] = 0;
        pixel_data[119][56] = 0;
        pixel_data[119][57] = 0;
        pixel_data[119][58] = 0;
        pixel_data[119][59] = 0;
        pixel_data[119][60] = 0;
        pixel_data[119][61] = 0;
        pixel_data[119][62] = 0;
        pixel_data[119][63] = 0;
        pixel_data[119][64] = 0;
        pixel_data[119][65] = 0;
        pixel_data[119][66] = 0;
        pixel_data[119][67] = 0;
        pixel_data[119][68] = 0;
        pixel_data[119][69] = 0;
        pixel_data[119][70] = 0;
        pixel_data[119][71] = 0;
        pixel_data[119][72] = 0;
        pixel_data[119][73] = 0;
        pixel_data[119][74] = 0;
        pixel_data[119][75] = 0;
        pixel_data[119][76] = 0;
        pixel_data[119][77] = 0;
        pixel_data[119][78] = 0;
        pixel_data[119][79] = 0;
        pixel_data[119][80] = 0;
        pixel_data[119][81] = 0;
        pixel_data[119][82] = 0;
        pixel_data[119][83] = 0;
        pixel_data[119][84] = 0;
        pixel_data[119][85] = 0;
        pixel_data[119][86] = 0;
        pixel_data[119][87] = 0;
        pixel_data[119][88] = 0;
        pixel_data[119][89] = 0;
        pixel_data[119][90] = 0;
        pixel_data[119][91] = 0;
        pixel_data[119][92] = 0;
        pixel_data[119][93] = 0;
        pixel_data[119][94] = 0;
        pixel_data[119][95] = 0;
        pixel_data[119][96] = 0;
        pixel_data[119][97] = 0;
        pixel_data[119][98] = 0;
        pixel_data[119][99] = 0;
        pixel_data[119][100] = 0;
        pixel_data[119][101] = 0;
        pixel_data[119][102] = 0;
        pixel_data[119][103] = 0;
        pixel_data[119][104] = 0;
        pixel_data[119][105] = 0;
        pixel_data[119][106] = 0;
        pixel_data[119][107] = 0;
        pixel_data[119][108] = 0;
        pixel_data[119][109] = 0;
        pixel_data[119][110] = 0;
        pixel_data[119][111] = 0;
        pixel_data[119][112] = 0;
        pixel_data[119][113] = 0;
        pixel_data[119][114] = 0;
        pixel_data[119][115] = 0;
        pixel_data[119][116] = 0;
        pixel_data[119][117] = 0;
        pixel_data[119][118] = 0;
        pixel_data[119][119] = 0;
        pixel_data[119][120] = 0;
        pixel_data[119][121] = 0;
        pixel_data[119][122] = 0;
        pixel_data[119][123] = 0;
        pixel_data[119][124] = 0;
        pixel_data[119][125] = 0;
        pixel_data[119][126] = 0;
        pixel_data[119][127] = 0;
        pixel_data[119][128] = 0;
        pixel_data[119][129] = 0;
        pixel_data[119][130] = 0;
        pixel_data[119][131] = 0;
        pixel_data[119][132] = 0;
        pixel_data[119][133] = 0;
        pixel_data[119][134] = 0;
        pixel_data[119][135] = 0;
        pixel_data[119][136] = 0;
        pixel_data[119][137] = 0;
        pixel_data[119][138] = 0;
        pixel_data[119][139] = 0;
        pixel_data[119][140] = 0;
        pixel_data[119][141] = 0;
        pixel_data[119][142] = 0;
        pixel_data[119][143] = 0;
        pixel_data[119][144] = 0;
        pixel_data[119][145] = 0;
        pixel_data[119][146] = 0;
        pixel_data[119][147] = 0;
        pixel_data[119][148] = 0;
        pixel_data[119][149] = 0;
        pixel_data[119][150] = 0;
        pixel_data[119][151] = 0;
        pixel_data[119][152] = 0;
        pixel_data[119][153] = 0;
        pixel_data[119][154] = 0;
        pixel_data[119][155] = 0;
        pixel_data[119][156] = 0;
        pixel_data[119][157] = 0;
        pixel_data[119][158] = 0;
        pixel_data[119][159] = 0;
        pixel_data[119][160] = 0;
        pixel_data[119][161] = 0;
        pixel_data[119][162] = 0;
        pixel_data[119][163] = 0;
        pixel_data[119][164] = 0;
        pixel_data[119][165] = 0;
        pixel_data[119][166] = 0;
        pixel_data[119][167] = 0;
        pixel_data[119][168] = 0;
        pixel_data[119][169] = 0;
        pixel_data[119][170] = 0;
        pixel_data[119][171] = 0;
        pixel_data[119][172] = 0;
        pixel_data[119][173] = 0;
        pixel_data[119][174] = 0;
        pixel_data[119][175] = 0;
        pixel_data[119][176] = 0;
        pixel_data[119][177] = 0;
        pixel_data[119][178] = 0;
        pixel_data[119][179] = 0;
        pixel_data[119][180] = 0;
        pixel_data[119][181] = 0;
        pixel_data[119][182] = 0;
        pixel_data[119][183] = 0;
        pixel_data[119][184] = 0;
        pixel_data[119][185] = 0;
        pixel_data[119][186] = 0;
        pixel_data[119][187] = 0;
        pixel_data[119][188] = 0;
        pixel_data[119][189] = 0;
        pixel_data[119][190] = 0;
        pixel_data[119][191] = 0;
        pixel_data[119][192] = 0;
        pixel_data[119][193] = 0;
        pixel_data[119][194] = 0;
        pixel_data[119][195] = 0;
        pixel_data[119][196] = 0;
        pixel_data[119][197] = 0;
        pixel_data[119][198] = 0;
        pixel_data[119][199] = 0; // y=119
        pixel_data[120][0] = 0;
        pixel_data[120][1] = 0;
        pixel_data[120][2] = 0;
        pixel_data[120][3] = 0;
        pixel_data[120][4] = 0;
        pixel_data[120][5] = 0;
        pixel_data[120][6] = 0;
        pixel_data[120][7] = 0;
        pixel_data[120][8] = 0;
        pixel_data[120][9] = 0;
        pixel_data[120][10] = 0;
        pixel_data[120][11] = 0;
        pixel_data[120][12] = 0;
        pixel_data[120][13] = 0;
        pixel_data[120][14] = 0;
        pixel_data[120][15] = 0;
        pixel_data[120][16] = 0;
        pixel_data[120][17] = 0;
        pixel_data[120][18] = 0;
        pixel_data[120][19] = 0;
        pixel_data[120][20] = 0;
        pixel_data[120][21] = 0;
        pixel_data[120][22] = 0;
        pixel_data[120][23] = 0;
        pixel_data[120][24] = 0;
        pixel_data[120][25] = 0;
        pixel_data[120][26] = 0;
        pixel_data[120][27] = 0;
        pixel_data[120][28] = 0;
        pixel_data[120][29] = 0;
        pixel_data[120][30] = 0;
        pixel_data[120][31] = 0;
        pixel_data[120][32] = 0;
        pixel_data[120][33] = 0;
        pixel_data[120][34] = 0;
        pixel_data[120][35] = 0;
        pixel_data[120][36] = 0;
        pixel_data[120][37] = 0;
        pixel_data[120][38] = 0;
        pixel_data[120][39] = 0;
        pixel_data[120][40] = 0;
        pixel_data[120][41] = 0;
        pixel_data[120][42] = 0;
        pixel_data[120][43] = 0;
        pixel_data[120][44] = 0;
        pixel_data[120][45] = 0;
        pixel_data[120][46] = 0;
        pixel_data[120][47] = 0;
        pixel_data[120][48] = 0;
        pixel_data[120][49] = 0;
        pixel_data[120][50] = 0;
        pixel_data[120][51] = 0;
        pixel_data[120][52] = 0;
        pixel_data[120][53] = 0;
        pixel_data[120][54] = 0;
        pixel_data[120][55] = 0;
        pixel_data[120][56] = 0;
        pixel_data[120][57] = 0;
        pixel_data[120][58] = 0;
        pixel_data[120][59] = 0;
        pixel_data[120][60] = 0;
        pixel_data[120][61] = 0;
        pixel_data[120][62] = 0;
        pixel_data[120][63] = 0;
        pixel_data[120][64] = 0;
        pixel_data[120][65] = 0;
        pixel_data[120][66] = 0;
        pixel_data[120][67] = 0;
        pixel_data[120][68] = 0;
        pixel_data[120][69] = 0;
        pixel_data[120][70] = 0;
        pixel_data[120][71] = 0;
        pixel_data[120][72] = 0;
        pixel_data[120][73] = 0;
        pixel_data[120][74] = 0;
        pixel_data[120][75] = 0;
        pixel_data[120][76] = 0;
        pixel_data[120][77] = 0;
        pixel_data[120][78] = 0;
        pixel_data[120][79] = 0;
        pixel_data[120][80] = 0;
        pixel_data[120][81] = 0;
        pixel_data[120][82] = 0;
        pixel_data[120][83] = 0;
        pixel_data[120][84] = 0;
        pixel_data[120][85] = 0;
        pixel_data[120][86] = 0;
        pixel_data[120][87] = 0;
        pixel_data[120][88] = 0;
        pixel_data[120][89] = 0;
        pixel_data[120][90] = 0;
        pixel_data[120][91] = 0;
        pixel_data[120][92] = 0;
        pixel_data[120][93] = 0;
        pixel_data[120][94] = 0;
        pixel_data[120][95] = 0;
        pixel_data[120][96] = 0;
        pixel_data[120][97] = 0;
        pixel_data[120][98] = 0;
        pixel_data[120][99] = 0;
        pixel_data[120][100] = 0;
        pixel_data[120][101] = 0;
        pixel_data[120][102] = 0;
        pixel_data[120][103] = 0;
        pixel_data[120][104] = 0;
        pixel_data[120][105] = 0;
        pixel_data[120][106] = 0;
        pixel_data[120][107] = 0;
        pixel_data[120][108] = 0;
        pixel_data[120][109] = 0;
        pixel_data[120][110] = 0;
        pixel_data[120][111] = 0;
        pixel_data[120][112] = 0;
        pixel_data[120][113] = 0;
        pixel_data[120][114] = 0;
        pixel_data[120][115] = 0;
        pixel_data[120][116] = 0;
        pixel_data[120][117] = 0;
        pixel_data[120][118] = 0;
        pixel_data[120][119] = 0;
        pixel_data[120][120] = 0;
        pixel_data[120][121] = 0;
        pixel_data[120][122] = 0;
        pixel_data[120][123] = 0;
        pixel_data[120][124] = 0;
        pixel_data[120][125] = 0;
        pixel_data[120][126] = 0;
        pixel_data[120][127] = 0;
        pixel_data[120][128] = 0;
        pixel_data[120][129] = 0;
        pixel_data[120][130] = 0;
        pixel_data[120][131] = 0;
        pixel_data[120][132] = 0;
        pixel_data[120][133] = 0;
        pixel_data[120][134] = 0;
        pixel_data[120][135] = 0;
        pixel_data[120][136] = 0;
        pixel_data[120][137] = 0;
        pixel_data[120][138] = 0;
        pixel_data[120][139] = 0;
        pixel_data[120][140] = 0;
        pixel_data[120][141] = 0;
        pixel_data[120][142] = 0;
        pixel_data[120][143] = 0;
        pixel_data[120][144] = 0;
        pixel_data[120][145] = 0;
        pixel_data[120][146] = 0;
        pixel_data[120][147] = 0;
        pixel_data[120][148] = 0;
        pixel_data[120][149] = 0;
        pixel_data[120][150] = 0;
        pixel_data[120][151] = 0;
        pixel_data[120][152] = 0;
        pixel_data[120][153] = 0;
        pixel_data[120][154] = 0;
        pixel_data[120][155] = 0;
        pixel_data[120][156] = 0;
        pixel_data[120][157] = 0;
        pixel_data[120][158] = 0;
        pixel_data[120][159] = 0;
        pixel_data[120][160] = 0;
        pixel_data[120][161] = 0;
        pixel_data[120][162] = 0;
        pixel_data[120][163] = 0;
        pixel_data[120][164] = 0;
        pixel_data[120][165] = 0;
        pixel_data[120][166] = 0;
        pixel_data[120][167] = 0;
        pixel_data[120][168] = 0;
        pixel_data[120][169] = 0;
        pixel_data[120][170] = 0;
        pixel_data[120][171] = 0;
        pixel_data[120][172] = 0;
        pixel_data[120][173] = 0;
        pixel_data[120][174] = 0;
        pixel_data[120][175] = 0;
        pixel_data[120][176] = 0;
        pixel_data[120][177] = 0;
        pixel_data[120][178] = 0;
        pixel_data[120][179] = 0;
        pixel_data[120][180] = 0;
        pixel_data[120][181] = 0;
        pixel_data[120][182] = 0;
        pixel_data[120][183] = 0;
        pixel_data[120][184] = 0;
        pixel_data[120][185] = 0;
        pixel_data[120][186] = 0;
        pixel_data[120][187] = 0;
        pixel_data[120][188] = 0;
        pixel_data[120][189] = 0;
        pixel_data[120][190] = 0;
        pixel_data[120][191] = 0;
        pixel_data[120][192] = 0;
        pixel_data[120][193] = 0;
        pixel_data[120][194] = 0;
        pixel_data[120][195] = 0;
        pixel_data[120][196] = 0;
        pixel_data[120][197] = 0;
        pixel_data[120][198] = 0;
        pixel_data[120][199] = 0; // y=120
        pixel_data[121][0] = 0;
        pixel_data[121][1] = 0;
        pixel_data[121][2] = 0;
        pixel_data[121][3] = 0;
        pixel_data[121][4] = 0;
        pixel_data[121][5] = 0;
        pixel_data[121][6] = 0;
        pixel_data[121][7] = 0;
        pixel_data[121][8] = 0;
        pixel_data[121][9] = 0;
        pixel_data[121][10] = 0;
        pixel_data[121][11] = 0;
        pixel_data[121][12] = 0;
        pixel_data[121][13] = 0;
        pixel_data[121][14] = 0;
        pixel_data[121][15] = 0;
        pixel_data[121][16] = 0;
        pixel_data[121][17] = 0;
        pixel_data[121][18] = 0;
        pixel_data[121][19] = 0;
        pixel_data[121][20] = 0;
        pixel_data[121][21] = 0;
        pixel_data[121][22] = 0;
        pixel_data[121][23] = 0;
        pixel_data[121][24] = 0;
        pixel_data[121][25] = 0;
        pixel_data[121][26] = 0;
        pixel_data[121][27] = 0;
        pixel_data[121][28] = 0;
        pixel_data[121][29] = 0;
        pixel_data[121][30] = 0;
        pixel_data[121][31] = 0;
        pixel_data[121][32] = 0;
        pixel_data[121][33] = 0;
        pixel_data[121][34] = 0;
        pixel_data[121][35] = 0;
        pixel_data[121][36] = 0;
        pixel_data[121][37] = 0;
        pixel_data[121][38] = 0;
        pixel_data[121][39] = 0;
        pixel_data[121][40] = 0;
        pixel_data[121][41] = 0;
        pixel_data[121][42] = 0;
        pixel_data[121][43] = 0;
        pixel_data[121][44] = 0;
        pixel_data[121][45] = 0;
        pixel_data[121][46] = 0;
        pixel_data[121][47] = 0;
        pixel_data[121][48] = 0;
        pixel_data[121][49] = 0;
        pixel_data[121][50] = 0;
        pixel_data[121][51] = 0;
        pixel_data[121][52] = 0;
        pixel_data[121][53] = 0;
        pixel_data[121][54] = 0;
        pixel_data[121][55] = 0;
        pixel_data[121][56] = 0;
        pixel_data[121][57] = 0;
        pixel_data[121][58] = 0;
        pixel_data[121][59] = 0;
        pixel_data[121][60] = 0;
        pixel_data[121][61] = 0;
        pixel_data[121][62] = 0;
        pixel_data[121][63] = 0;
        pixel_data[121][64] = 0;
        pixel_data[121][65] = 0;
        pixel_data[121][66] = 0;
        pixel_data[121][67] = 0;
        pixel_data[121][68] = 0;
        pixel_data[121][69] = 0;
        pixel_data[121][70] = 0;
        pixel_data[121][71] = 0;
        pixel_data[121][72] = 0;
        pixel_data[121][73] = 0;
        pixel_data[121][74] = 0;
        pixel_data[121][75] = 0;
        pixel_data[121][76] = 0;
        pixel_data[121][77] = 0;
        pixel_data[121][78] = 0;
        pixel_data[121][79] = 0;
        pixel_data[121][80] = 0;
        pixel_data[121][81] = 0;
        pixel_data[121][82] = 0;
        pixel_data[121][83] = 0;
        pixel_data[121][84] = 0;
        pixel_data[121][85] = 0;
        pixel_data[121][86] = 0;
        pixel_data[121][87] = 0;
        pixel_data[121][88] = 0;
        pixel_data[121][89] = 0;
        pixel_data[121][90] = 0;
        pixel_data[121][91] = 0;
        pixel_data[121][92] = 0;
        pixel_data[121][93] = 0;
        pixel_data[121][94] = 0;
        pixel_data[121][95] = 0;
        pixel_data[121][96] = 0;
        pixel_data[121][97] = 0;
        pixel_data[121][98] = 0;
        pixel_data[121][99] = 0;
        pixel_data[121][100] = 0;
        pixel_data[121][101] = 0;
        pixel_data[121][102] = 0;
        pixel_data[121][103] = 0;
        pixel_data[121][104] = 0;
        pixel_data[121][105] = 0;
        pixel_data[121][106] = 0;
        pixel_data[121][107] = 0;
        pixel_data[121][108] = 0;
        pixel_data[121][109] = 0;
        pixel_data[121][110] = 0;
        pixel_data[121][111] = 0;
        pixel_data[121][112] = 0;
        pixel_data[121][113] = 0;
        pixel_data[121][114] = 0;
        pixel_data[121][115] = 0;
        pixel_data[121][116] = 0;
        pixel_data[121][117] = 0;
        pixel_data[121][118] = 0;
        pixel_data[121][119] = 0;
        pixel_data[121][120] = 0;
        pixel_data[121][121] = 0;
        pixel_data[121][122] = 0;
        pixel_data[121][123] = 0;
        pixel_data[121][124] = 0;
        pixel_data[121][125] = 0;
        pixel_data[121][126] = 0;
        pixel_data[121][127] = 0;
        pixel_data[121][128] = 0;
        pixel_data[121][129] = 0;
        pixel_data[121][130] = 0;
        pixel_data[121][131] = 0;
        pixel_data[121][132] = 0;
        pixel_data[121][133] = 0;
        pixel_data[121][134] = 0;
        pixel_data[121][135] = 0;
        pixel_data[121][136] = 0;
        pixel_data[121][137] = 0;
        pixel_data[121][138] = 0;
        pixel_data[121][139] = 0;
        pixel_data[121][140] = 0;
        pixel_data[121][141] = 0;
        pixel_data[121][142] = 0;
        pixel_data[121][143] = 0;
        pixel_data[121][144] = 0;
        pixel_data[121][145] = 0;
        pixel_data[121][146] = 0;
        pixel_data[121][147] = 0;
        pixel_data[121][148] = 0;
        pixel_data[121][149] = 0;
        pixel_data[121][150] = 0;
        pixel_data[121][151] = 0;
        pixel_data[121][152] = 0;
        pixel_data[121][153] = 0;
        pixel_data[121][154] = 0;
        pixel_data[121][155] = 0;
        pixel_data[121][156] = 0;
        pixel_data[121][157] = 0;
        pixel_data[121][158] = 0;
        pixel_data[121][159] = 0;
        pixel_data[121][160] = 0;
        pixel_data[121][161] = 0;
        pixel_data[121][162] = 0;
        pixel_data[121][163] = 0;
        pixel_data[121][164] = 0;
        pixel_data[121][165] = 0;
        pixel_data[121][166] = 0;
        pixel_data[121][167] = 0;
        pixel_data[121][168] = 0;
        pixel_data[121][169] = 0;
        pixel_data[121][170] = 0;
        pixel_data[121][171] = 0;
        pixel_data[121][172] = 0;
        pixel_data[121][173] = 0;
        pixel_data[121][174] = 0;
        pixel_data[121][175] = 0;
        pixel_data[121][176] = 0;
        pixel_data[121][177] = 0;
        pixel_data[121][178] = 0;
        pixel_data[121][179] = 0;
        pixel_data[121][180] = 0;
        pixel_data[121][181] = 0;
        pixel_data[121][182] = 0;
        pixel_data[121][183] = 0;
        pixel_data[121][184] = 0;
        pixel_data[121][185] = 0;
        pixel_data[121][186] = 0;
        pixel_data[121][187] = 0;
        pixel_data[121][188] = 0;
        pixel_data[121][189] = 0;
        pixel_data[121][190] = 0;
        pixel_data[121][191] = 0;
        pixel_data[121][192] = 0;
        pixel_data[121][193] = 0;
        pixel_data[121][194] = 0;
        pixel_data[121][195] = 0;
        pixel_data[121][196] = 0;
        pixel_data[121][197] = 0;
        pixel_data[121][198] = 0;
        pixel_data[121][199] = 0; // y=121
        pixel_data[122][0] = 0;
        pixel_data[122][1] = 0;
        pixel_data[122][2] = 0;
        pixel_data[122][3] = 0;
        pixel_data[122][4] = 0;
        pixel_data[122][5] = 0;
        pixel_data[122][6] = 0;
        pixel_data[122][7] = 0;
        pixel_data[122][8] = 0;
        pixel_data[122][9] = 0;
        pixel_data[122][10] = 0;
        pixel_data[122][11] = 0;
        pixel_data[122][12] = 0;
        pixel_data[122][13] = 0;
        pixel_data[122][14] = 0;
        pixel_data[122][15] = 0;
        pixel_data[122][16] = 0;
        pixel_data[122][17] = 0;
        pixel_data[122][18] = 0;
        pixel_data[122][19] = 0;
        pixel_data[122][20] = 0;
        pixel_data[122][21] = 0;
        pixel_data[122][22] = 0;
        pixel_data[122][23] = 0;
        pixel_data[122][24] = 0;
        pixel_data[122][25] = 0;
        pixel_data[122][26] = 0;
        pixel_data[122][27] = 0;
        pixel_data[122][28] = 0;
        pixel_data[122][29] = 0;
        pixel_data[122][30] = 0;
        pixel_data[122][31] = 0;
        pixel_data[122][32] = 0;
        pixel_data[122][33] = 0;
        pixel_data[122][34] = 0;
        pixel_data[122][35] = 0;
        pixel_data[122][36] = 0;
        pixel_data[122][37] = 0;
        pixel_data[122][38] = 0;
        pixel_data[122][39] = 0;
        pixel_data[122][40] = 0;
        pixel_data[122][41] = 0;
        pixel_data[122][42] = 0;
        pixel_data[122][43] = 0;
        pixel_data[122][44] = 0;
        pixel_data[122][45] = 0;
        pixel_data[122][46] = 0;
        pixel_data[122][47] = 0;
        pixel_data[122][48] = 0;
        pixel_data[122][49] = 0;
        pixel_data[122][50] = 0;
        pixel_data[122][51] = 0;
        pixel_data[122][52] = 0;
        pixel_data[122][53] = 0;
        pixel_data[122][54] = 0;
        pixel_data[122][55] = 0;
        pixel_data[122][56] = 0;
        pixel_data[122][57] = 0;
        pixel_data[122][58] = 0;
        pixel_data[122][59] = 0;
        pixel_data[122][60] = 0;
        pixel_data[122][61] = 0;
        pixel_data[122][62] = 0;
        pixel_data[122][63] = 0;
        pixel_data[122][64] = 0;
        pixel_data[122][65] = 0;
        pixel_data[122][66] = 0;
        pixel_data[122][67] = 0;
        pixel_data[122][68] = 0;
        pixel_data[122][69] = 0;
        pixel_data[122][70] = 0;
        pixel_data[122][71] = 0;
        pixel_data[122][72] = 0;
        pixel_data[122][73] = 0;
        pixel_data[122][74] = 0;
        pixel_data[122][75] = 0;
        pixel_data[122][76] = 0;
        pixel_data[122][77] = 0;
        pixel_data[122][78] = 0;
        pixel_data[122][79] = 0;
        pixel_data[122][80] = 0;
        pixel_data[122][81] = 0;
        pixel_data[122][82] = 0;
        pixel_data[122][83] = 0;
        pixel_data[122][84] = 0;
        pixel_data[122][85] = 0;
        pixel_data[122][86] = 0;
        pixel_data[122][87] = 0;
        pixel_data[122][88] = 0;
        pixel_data[122][89] = 0;
        pixel_data[122][90] = 0;
        pixel_data[122][91] = 0;
        pixel_data[122][92] = 0;
        pixel_data[122][93] = 0;
        pixel_data[122][94] = 0;
        pixel_data[122][95] = 0;
        pixel_data[122][96] = 0;
        pixel_data[122][97] = 0;
        pixel_data[122][98] = 0;
        pixel_data[122][99] = 0;
        pixel_data[122][100] = 0;
        pixel_data[122][101] = 0;
        pixel_data[122][102] = 0;
        pixel_data[122][103] = 0;
        pixel_data[122][104] = 0;
        pixel_data[122][105] = 0;
        pixel_data[122][106] = 0;
        pixel_data[122][107] = 0;
        pixel_data[122][108] = 0;
        pixel_data[122][109] = 0;
        pixel_data[122][110] = 0;
        pixel_data[122][111] = 0;
        pixel_data[122][112] = 0;
        pixel_data[122][113] = 0;
        pixel_data[122][114] = 0;
        pixel_data[122][115] = 0;
        pixel_data[122][116] = 0;
        pixel_data[122][117] = 0;
        pixel_data[122][118] = 0;
        pixel_data[122][119] = 0;
        pixel_data[122][120] = 0;
        pixel_data[122][121] = 0;
        pixel_data[122][122] = 0;
        pixel_data[122][123] = 0;
        pixel_data[122][124] = 0;
        pixel_data[122][125] = 0;
        pixel_data[122][126] = 0;
        pixel_data[122][127] = 0;
        pixel_data[122][128] = 0;
        pixel_data[122][129] = 0;
        pixel_data[122][130] = 0;
        pixel_data[122][131] = 0;
        pixel_data[122][132] = 0;
        pixel_data[122][133] = 0;
        pixel_data[122][134] = 0;
        pixel_data[122][135] = 0;
        pixel_data[122][136] = 0;
        pixel_data[122][137] = 0;
        pixel_data[122][138] = 0;
        pixel_data[122][139] = 0;
        pixel_data[122][140] = 0;
        pixel_data[122][141] = 0;
        pixel_data[122][142] = 0;
        pixel_data[122][143] = 0;
        pixel_data[122][144] = 0;
        pixel_data[122][145] = 0;
        pixel_data[122][146] = 0;
        pixel_data[122][147] = 0;
        pixel_data[122][148] = 0;
        pixel_data[122][149] = 0;
        pixel_data[122][150] = 0;
        pixel_data[122][151] = 0;
        pixel_data[122][152] = 0;
        pixel_data[122][153] = 0;
        pixel_data[122][154] = 0;
        pixel_data[122][155] = 0;
        pixel_data[122][156] = 0;
        pixel_data[122][157] = 0;
        pixel_data[122][158] = 0;
        pixel_data[122][159] = 0;
        pixel_data[122][160] = 0;
        pixel_data[122][161] = 0;
        pixel_data[122][162] = 0;
        pixel_data[122][163] = 0;
        pixel_data[122][164] = 0;
        pixel_data[122][165] = 0;
        pixel_data[122][166] = 0;
        pixel_data[122][167] = 0;
        pixel_data[122][168] = 0;
        pixel_data[122][169] = 0;
        pixel_data[122][170] = 0;
        pixel_data[122][171] = 0;
        pixel_data[122][172] = 0;
        pixel_data[122][173] = 0;
        pixel_data[122][174] = 0;
        pixel_data[122][175] = 0;
        pixel_data[122][176] = 0;
        pixel_data[122][177] = 0;
        pixel_data[122][178] = 0;
        pixel_data[122][179] = 0;
        pixel_data[122][180] = 0;
        pixel_data[122][181] = 0;
        pixel_data[122][182] = 0;
        pixel_data[122][183] = 0;
        pixel_data[122][184] = 0;
        pixel_data[122][185] = 0;
        pixel_data[122][186] = 0;
        pixel_data[122][187] = 0;
        pixel_data[122][188] = 0;
        pixel_data[122][189] = 0;
        pixel_data[122][190] = 0;
        pixel_data[122][191] = 0;
        pixel_data[122][192] = 0;
        pixel_data[122][193] = 0;
        pixel_data[122][194] = 0;
        pixel_data[122][195] = 0;
        pixel_data[122][196] = 0;
        pixel_data[122][197] = 0;
        pixel_data[122][198] = 0;
        pixel_data[122][199] = 0; // y=122
        pixel_data[123][0] = 0;
        pixel_data[123][1] = 0;
        pixel_data[123][2] = 0;
        pixel_data[123][3] = 0;
        pixel_data[123][4] = 0;
        pixel_data[123][5] = 0;
        pixel_data[123][6] = 0;
        pixel_data[123][7] = 0;
        pixel_data[123][8] = 0;
        pixel_data[123][9] = 0;
        pixel_data[123][10] = 0;
        pixel_data[123][11] = 0;
        pixel_data[123][12] = 0;
        pixel_data[123][13] = 0;
        pixel_data[123][14] = 0;
        pixel_data[123][15] = 0;
        pixel_data[123][16] = 0;
        pixel_data[123][17] = 0;
        pixel_data[123][18] = 0;
        pixel_data[123][19] = 0;
        pixel_data[123][20] = 0;
        pixel_data[123][21] = 0;
        pixel_data[123][22] = 0;
        pixel_data[123][23] = 0;
        pixel_data[123][24] = 0;
        pixel_data[123][25] = 0;
        pixel_data[123][26] = 0;
        pixel_data[123][27] = 0;
        pixel_data[123][28] = 0;
        pixel_data[123][29] = 0;
        pixel_data[123][30] = 0;
        pixel_data[123][31] = 0;
        pixel_data[123][32] = 0;
        pixel_data[123][33] = 0;
        pixel_data[123][34] = 0;
        pixel_data[123][35] = 0;
        pixel_data[123][36] = 0;
        pixel_data[123][37] = 0;
        pixel_data[123][38] = 0;
        pixel_data[123][39] = 0;
        pixel_data[123][40] = 0;
        pixel_data[123][41] = 0;
        pixel_data[123][42] = 0;
        pixel_data[123][43] = 0;
        pixel_data[123][44] = 0;
        pixel_data[123][45] = 0;
        pixel_data[123][46] = 0;
        pixel_data[123][47] = 0;
        pixel_data[123][48] = 0;
        pixel_data[123][49] = 0;
        pixel_data[123][50] = 0;
        pixel_data[123][51] = 0;
        pixel_data[123][52] = 0;
        pixel_data[123][53] = 0;
        pixel_data[123][54] = 0;
        pixel_data[123][55] = 0;
        pixel_data[123][56] = 0;
        pixel_data[123][57] = 0;
        pixel_data[123][58] = 0;
        pixel_data[123][59] = 0;
        pixel_data[123][60] = 0;
        pixel_data[123][61] = 0;
        pixel_data[123][62] = 0;
        pixel_data[123][63] = 0;
        pixel_data[123][64] = 0;
        pixel_data[123][65] = 0;
        pixel_data[123][66] = 0;
        pixel_data[123][67] = 0;
        pixel_data[123][68] = 0;
        pixel_data[123][69] = 0;
        pixel_data[123][70] = 0;
        pixel_data[123][71] = 0;
        pixel_data[123][72] = 0;
        pixel_data[123][73] = 0;
        pixel_data[123][74] = 0;
        pixel_data[123][75] = 0;
        pixel_data[123][76] = 0;
        pixel_data[123][77] = 0;
        pixel_data[123][78] = 0;
        pixel_data[123][79] = 0;
        pixel_data[123][80] = 0;
        pixel_data[123][81] = 0;
        pixel_data[123][82] = 0;
        pixel_data[123][83] = 0;
        pixel_data[123][84] = 0;
        pixel_data[123][85] = 0;
        pixel_data[123][86] = 0;
        pixel_data[123][87] = 0;
        pixel_data[123][88] = 0;
        pixel_data[123][89] = 0;
        pixel_data[123][90] = 0;
        pixel_data[123][91] = 0;
        pixel_data[123][92] = 0;
        pixel_data[123][93] = 0;
        pixel_data[123][94] = 0;
        pixel_data[123][95] = 0;
        pixel_data[123][96] = 0;
        pixel_data[123][97] = 0;
        pixel_data[123][98] = 0;
        pixel_data[123][99] = 0;
        pixel_data[123][100] = 0;
        pixel_data[123][101] = 0;
        pixel_data[123][102] = 0;
        pixel_data[123][103] = 0;
        pixel_data[123][104] = 0;
        pixel_data[123][105] = 0;
        pixel_data[123][106] = 0;
        pixel_data[123][107] = 0;
        pixel_data[123][108] = 0;
        pixel_data[123][109] = 0;
        pixel_data[123][110] = 0;
        pixel_data[123][111] = 0;
        pixel_data[123][112] = 0;
        pixel_data[123][113] = 0;
        pixel_data[123][114] = 0;
        pixel_data[123][115] = 0;
        pixel_data[123][116] = 0;
        pixel_data[123][117] = 0;
        pixel_data[123][118] = 0;
        pixel_data[123][119] = 0;
        pixel_data[123][120] = 0;
        pixel_data[123][121] = 0;
        pixel_data[123][122] = 0;
        pixel_data[123][123] = 0;
        pixel_data[123][124] = 0;
        pixel_data[123][125] = 0;
        pixel_data[123][126] = 0;
        pixel_data[123][127] = 0;
        pixel_data[123][128] = 0;
        pixel_data[123][129] = 0;
        pixel_data[123][130] = 0;
        pixel_data[123][131] = 0;
        pixel_data[123][132] = 0;
        pixel_data[123][133] = 0;
        pixel_data[123][134] = 0;
        pixel_data[123][135] = 0;
        pixel_data[123][136] = 0;
        pixel_data[123][137] = 0;
        pixel_data[123][138] = 0;
        pixel_data[123][139] = 0;
        pixel_data[123][140] = 0;
        pixel_data[123][141] = 0;
        pixel_data[123][142] = 0;
        pixel_data[123][143] = 0;
        pixel_data[123][144] = 0;
        pixel_data[123][145] = 0;
        pixel_data[123][146] = 0;
        pixel_data[123][147] = 0;
        pixel_data[123][148] = 0;
        pixel_data[123][149] = 0;
        pixel_data[123][150] = 0;
        pixel_data[123][151] = 0;
        pixel_data[123][152] = 0;
        pixel_data[123][153] = 0;
        pixel_data[123][154] = 0;
        pixel_data[123][155] = 0;
        pixel_data[123][156] = 0;
        pixel_data[123][157] = 0;
        pixel_data[123][158] = 0;
        pixel_data[123][159] = 0;
        pixel_data[123][160] = 0;
        pixel_data[123][161] = 0;
        pixel_data[123][162] = 0;
        pixel_data[123][163] = 0;
        pixel_data[123][164] = 0;
        pixel_data[123][165] = 0;
        pixel_data[123][166] = 0;
        pixel_data[123][167] = 0;
        pixel_data[123][168] = 0;
        pixel_data[123][169] = 0;
        pixel_data[123][170] = 0;
        pixel_data[123][171] = 0;
        pixel_data[123][172] = 0;
        pixel_data[123][173] = 0;
        pixel_data[123][174] = 0;
        pixel_data[123][175] = 0;
        pixel_data[123][176] = 0;
        pixel_data[123][177] = 0;
        pixel_data[123][178] = 0;
        pixel_data[123][179] = 0;
        pixel_data[123][180] = 0;
        pixel_data[123][181] = 0;
        pixel_data[123][182] = 0;
        pixel_data[123][183] = 0;
        pixel_data[123][184] = 0;
        pixel_data[123][185] = 0;
        pixel_data[123][186] = 0;
        pixel_data[123][187] = 0;
        pixel_data[123][188] = 0;
        pixel_data[123][189] = 0;
        pixel_data[123][190] = 0;
        pixel_data[123][191] = 0;
        pixel_data[123][192] = 0;
        pixel_data[123][193] = 0;
        pixel_data[123][194] = 0;
        pixel_data[123][195] = 0;
        pixel_data[123][196] = 0;
        pixel_data[123][197] = 0;
        pixel_data[123][198] = 0;
        pixel_data[123][199] = 0; // y=123
        pixel_data[124][0] = 0;
        pixel_data[124][1] = 0;
        pixel_data[124][2] = 0;
        pixel_data[124][3] = 0;
        pixel_data[124][4] = 0;
        pixel_data[124][5] = 0;
        pixel_data[124][6] = 0;
        pixel_data[124][7] = 0;
        pixel_data[124][8] = 0;
        pixel_data[124][9] = 0;
        pixel_data[124][10] = 0;
        pixel_data[124][11] = 0;
        pixel_data[124][12] = 0;
        pixel_data[124][13] = 0;
        pixel_data[124][14] = 0;
        pixel_data[124][15] = 0;
        pixel_data[124][16] = 0;
        pixel_data[124][17] = 0;
        pixel_data[124][18] = 0;
        pixel_data[124][19] = 0;
        pixel_data[124][20] = 0;
        pixel_data[124][21] = 0;
        pixel_data[124][22] = 0;
        pixel_data[124][23] = 0;
        pixel_data[124][24] = 0;
        pixel_data[124][25] = 0;
        pixel_data[124][26] = 0;
        pixel_data[124][27] = 0;
        pixel_data[124][28] = 0;
        pixel_data[124][29] = 0;
        pixel_data[124][30] = 0;
        pixel_data[124][31] = 0;
        pixel_data[124][32] = 0;
        pixel_data[124][33] = 0;
        pixel_data[124][34] = 0;
        pixel_data[124][35] = 0;
        pixel_data[124][36] = 0;
        pixel_data[124][37] = 0;
        pixel_data[124][38] = 0;
        pixel_data[124][39] = 0;
        pixel_data[124][40] = 0;
        pixel_data[124][41] = 0;
        pixel_data[124][42] = 0;
        pixel_data[124][43] = 0;
        pixel_data[124][44] = 0;
        pixel_data[124][45] = 0;
        pixel_data[124][46] = 0;
        pixel_data[124][47] = 0;
        pixel_data[124][48] = 0;
        pixel_data[124][49] = 0;
        pixel_data[124][50] = 0;
        pixel_data[124][51] = 0;
        pixel_data[124][52] = 0;
        pixel_data[124][53] = 0;
        pixel_data[124][54] = 0;
        pixel_data[124][55] = 0;
        pixel_data[124][56] = 0;
        pixel_data[124][57] = 0;
        pixel_data[124][58] = 0;
        pixel_data[124][59] = 0;
        pixel_data[124][60] = 0;
        pixel_data[124][61] = 0;
        pixel_data[124][62] = 0;
        pixel_data[124][63] = 0;
        pixel_data[124][64] = 0;
        pixel_data[124][65] = 0;
        pixel_data[124][66] = 0;
        pixel_data[124][67] = 0;
        pixel_data[124][68] = 0;
        pixel_data[124][69] = 0;
        pixel_data[124][70] = 0;
        pixel_data[124][71] = 0;
        pixel_data[124][72] = 0;
        pixel_data[124][73] = 0;
        pixel_data[124][74] = 0;
        pixel_data[124][75] = 0;
        pixel_data[124][76] = 0;
        pixel_data[124][77] = 0;
        pixel_data[124][78] = 0;
        pixel_data[124][79] = 0;
        pixel_data[124][80] = 0;
        pixel_data[124][81] = 0;
        pixel_data[124][82] = 0;
        pixel_data[124][83] = 0;
        pixel_data[124][84] = 0;
        pixel_data[124][85] = 0;
        pixel_data[124][86] = 0;
        pixel_data[124][87] = 0;
        pixel_data[124][88] = 0;
        pixel_data[124][89] = 0;
        pixel_data[124][90] = 0;
        pixel_data[124][91] = 0;
        pixel_data[124][92] = 0;
        pixel_data[124][93] = 0;
        pixel_data[124][94] = 0;
        pixel_data[124][95] = 0;
        pixel_data[124][96] = 0;
        pixel_data[124][97] = 0;
        pixel_data[124][98] = 0;
        pixel_data[124][99] = 0;
        pixel_data[124][100] = 0;
        pixel_data[124][101] = 0;
        pixel_data[124][102] = 0;
        pixel_data[124][103] = 0;
        pixel_data[124][104] = 0;
        pixel_data[124][105] = 0;
        pixel_data[124][106] = 0;
        pixel_data[124][107] = 0;
        pixel_data[124][108] = 0;
        pixel_data[124][109] = 0;
        pixel_data[124][110] = 0;
        pixel_data[124][111] = 0;
        pixel_data[124][112] = 0;
        pixel_data[124][113] = 0;
        pixel_data[124][114] = 0;
        pixel_data[124][115] = 0;
        pixel_data[124][116] = 0;
        pixel_data[124][117] = 0;
        pixel_data[124][118] = 0;
        pixel_data[124][119] = 0;
        pixel_data[124][120] = 0;
        pixel_data[124][121] = 0;
        pixel_data[124][122] = 0;
        pixel_data[124][123] = 0;
        pixel_data[124][124] = 0;
        pixel_data[124][125] = 0;
        pixel_data[124][126] = 0;
        pixel_data[124][127] = 0;
        pixel_data[124][128] = 0;
        pixel_data[124][129] = 0;
        pixel_data[124][130] = 0;
        pixel_data[124][131] = 0;
        pixel_data[124][132] = 0;
        pixel_data[124][133] = 0;
        pixel_data[124][134] = 0;
        pixel_data[124][135] = 0;
        pixel_data[124][136] = 0;
        pixel_data[124][137] = 0;
        pixel_data[124][138] = 0;
        pixel_data[124][139] = 0;
        pixel_data[124][140] = 0;
        pixel_data[124][141] = 0;
        pixel_data[124][142] = 0;
        pixel_data[124][143] = 0;
        pixel_data[124][144] = 0;
        pixel_data[124][145] = 0;
        pixel_data[124][146] = 0;
        pixel_data[124][147] = 0;
        pixel_data[124][148] = 0;
        pixel_data[124][149] = 0;
        pixel_data[124][150] = 0;
        pixel_data[124][151] = 0;
        pixel_data[124][152] = 0;
        pixel_data[124][153] = 0;
        pixel_data[124][154] = 0;
        pixel_data[124][155] = 0;
        pixel_data[124][156] = 0;
        pixel_data[124][157] = 0;
        pixel_data[124][158] = 0;
        pixel_data[124][159] = 0;
        pixel_data[124][160] = 0;
        pixel_data[124][161] = 0;
        pixel_data[124][162] = 0;
        pixel_data[124][163] = 0;
        pixel_data[124][164] = 0;
        pixel_data[124][165] = 0;
        pixel_data[124][166] = 0;
        pixel_data[124][167] = 0;
        pixel_data[124][168] = 0;
        pixel_data[124][169] = 0;
        pixel_data[124][170] = 0;
        pixel_data[124][171] = 0;
        pixel_data[124][172] = 0;
        pixel_data[124][173] = 0;
        pixel_data[124][174] = 0;
        pixel_data[124][175] = 0;
        pixel_data[124][176] = 0;
        pixel_data[124][177] = 0;
        pixel_data[124][178] = 0;
        pixel_data[124][179] = 0;
        pixel_data[124][180] = 0;
        pixel_data[124][181] = 0;
        pixel_data[124][182] = 0;
        pixel_data[124][183] = 0;
        pixel_data[124][184] = 0;
        pixel_data[124][185] = 0;
        pixel_data[124][186] = 0;
        pixel_data[124][187] = 0;
        pixel_data[124][188] = 0;
        pixel_data[124][189] = 0;
        pixel_data[124][190] = 0;
        pixel_data[124][191] = 0;
        pixel_data[124][192] = 0;
        pixel_data[124][193] = 0;
        pixel_data[124][194] = 0;
        pixel_data[124][195] = 0;
        pixel_data[124][196] = 0;
        pixel_data[124][197] = 0;
        pixel_data[124][198] = 0;
        pixel_data[124][199] = 0; // y=124
        pixel_data[125][0] = 0;
        pixel_data[125][1] = 0;
        pixel_data[125][2] = 0;
        pixel_data[125][3] = 0;
        pixel_data[125][4] = 0;
        pixel_data[125][5] = 0;
        pixel_data[125][6] = 0;
        pixel_data[125][7] = 0;
        pixel_data[125][8] = 0;
        pixel_data[125][9] = 0;
        pixel_data[125][10] = 0;
        pixel_data[125][11] = 0;
        pixel_data[125][12] = 0;
        pixel_data[125][13] = 0;
        pixel_data[125][14] = 0;
        pixel_data[125][15] = 0;
        pixel_data[125][16] = 0;
        pixel_data[125][17] = 0;
        pixel_data[125][18] = 0;
        pixel_data[125][19] = 0;
        pixel_data[125][20] = 0;
        pixel_data[125][21] = 0;
        pixel_data[125][22] = 0;
        pixel_data[125][23] = 0;
        pixel_data[125][24] = 0;
        pixel_data[125][25] = 0;
        pixel_data[125][26] = 0;
        pixel_data[125][27] = 0;
        pixel_data[125][28] = 0;
        pixel_data[125][29] = 0;
        pixel_data[125][30] = 0;
        pixel_data[125][31] = 0;
        pixel_data[125][32] = 0;
        pixel_data[125][33] = 0;
        pixel_data[125][34] = 0;
        pixel_data[125][35] = 0;
        pixel_data[125][36] = 0;
        pixel_data[125][37] = 0;
        pixel_data[125][38] = 0;
        pixel_data[125][39] = 0;
        pixel_data[125][40] = 0;
        pixel_data[125][41] = 0;
        pixel_data[125][42] = 0;
        pixel_data[125][43] = 0;
        pixel_data[125][44] = 0;
        pixel_data[125][45] = 0;
        pixel_data[125][46] = 0;
        pixel_data[125][47] = 0;
        pixel_data[125][48] = 0;
        pixel_data[125][49] = 0;
        pixel_data[125][50] = 0;
        pixel_data[125][51] = 0;
        pixel_data[125][52] = 0;
        pixel_data[125][53] = 0;
        pixel_data[125][54] = 0;
        pixel_data[125][55] = 0;
        pixel_data[125][56] = 0;
        pixel_data[125][57] = 0;
        pixel_data[125][58] = 0;
        pixel_data[125][59] = 0;
        pixel_data[125][60] = 0;
        pixel_data[125][61] = 0;
        pixel_data[125][62] = 0;
        pixel_data[125][63] = 0;
        pixel_data[125][64] = 0;
        pixel_data[125][65] = 0;
        pixel_data[125][66] = 0;
        pixel_data[125][67] = 0;
        pixel_data[125][68] = 0;
        pixel_data[125][69] = 0;
        pixel_data[125][70] = 0;
        pixel_data[125][71] = 0;
        pixel_data[125][72] = 0;
        pixel_data[125][73] = 0;
        pixel_data[125][74] = 0;
        pixel_data[125][75] = 0;
        pixel_data[125][76] = 0;
        pixel_data[125][77] = 0;
        pixel_data[125][78] = 0;
        pixel_data[125][79] = 0;
        pixel_data[125][80] = 0;
        pixel_data[125][81] = 0;
        pixel_data[125][82] = 0;
        pixel_data[125][83] = 0;
        pixel_data[125][84] = 0;
        pixel_data[125][85] = 0;
        pixel_data[125][86] = 0;
        pixel_data[125][87] = 0;
        pixel_data[125][88] = 0;
        pixel_data[125][89] = 0;
        pixel_data[125][90] = 0;
        pixel_data[125][91] = 0;
        pixel_data[125][92] = 0;
        pixel_data[125][93] = 0;
        pixel_data[125][94] = 0;
        pixel_data[125][95] = 0;
        pixel_data[125][96] = 0;
        pixel_data[125][97] = 0;
        pixel_data[125][98] = 0;
        pixel_data[125][99] = 0;
        pixel_data[125][100] = 0;
        pixel_data[125][101] = 0;
        pixel_data[125][102] = 0;
        pixel_data[125][103] = 0;
        pixel_data[125][104] = 0;
        pixel_data[125][105] = 0;
        pixel_data[125][106] = 0;
        pixel_data[125][107] = 0;
        pixel_data[125][108] = 0;
        pixel_data[125][109] = 0;
        pixel_data[125][110] = 0;
        pixel_data[125][111] = 0;
        pixel_data[125][112] = 0;
        pixel_data[125][113] = 0;
        pixel_data[125][114] = 0;
        pixel_data[125][115] = 0;
        pixel_data[125][116] = 0;
        pixel_data[125][117] = 0;
        pixel_data[125][118] = 0;
        pixel_data[125][119] = 0;
        pixel_data[125][120] = 0;
        pixel_data[125][121] = 0;
        pixel_data[125][122] = 0;
        pixel_data[125][123] = 0;
        pixel_data[125][124] = 0;
        pixel_data[125][125] = 0;
        pixel_data[125][126] = 0;
        pixel_data[125][127] = 0;
        pixel_data[125][128] = 0;
        pixel_data[125][129] = 0;
        pixel_data[125][130] = 0;
        pixel_data[125][131] = 0;
        pixel_data[125][132] = 0;
        pixel_data[125][133] = 0;
        pixel_data[125][134] = 0;
        pixel_data[125][135] = 0;
        pixel_data[125][136] = 0;
        pixel_data[125][137] = 0;
        pixel_data[125][138] = 0;
        pixel_data[125][139] = 0;
        pixel_data[125][140] = 0;
        pixel_data[125][141] = 0;
        pixel_data[125][142] = 0;
        pixel_data[125][143] = 0;
        pixel_data[125][144] = 0;
        pixel_data[125][145] = 0;
        pixel_data[125][146] = 0;
        pixel_data[125][147] = 0;
        pixel_data[125][148] = 0;
        pixel_data[125][149] = 0;
        pixel_data[125][150] = 0;
        pixel_data[125][151] = 0;
        pixel_data[125][152] = 0;
        pixel_data[125][153] = 0;
        pixel_data[125][154] = 0;
        pixel_data[125][155] = 0;
        pixel_data[125][156] = 0;
        pixel_data[125][157] = 0;
        pixel_data[125][158] = 0;
        pixel_data[125][159] = 0;
        pixel_data[125][160] = 0;
        pixel_data[125][161] = 0;
        pixel_data[125][162] = 0;
        pixel_data[125][163] = 0;
        pixel_data[125][164] = 0;
        pixel_data[125][165] = 0;
        pixel_data[125][166] = 0;
        pixel_data[125][167] = 0;
        pixel_data[125][168] = 0;
        pixel_data[125][169] = 0;
        pixel_data[125][170] = 0;
        pixel_data[125][171] = 0;
        pixel_data[125][172] = 0;
        pixel_data[125][173] = 0;
        pixel_data[125][174] = 0;
        pixel_data[125][175] = 0;
        pixel_data[125][176] = 0;
        pixel_data[125][177] = 0;
        pixel_data[125][178] = 0;
        pixel_data[125][179] = 0;
        pixel_data[125][180] = 0;
        pixel_data[125][181] = 0;
        pixel_data[125][182] = 0;
        pixel_data[125][183] = 0;
        pixel_data[125][184] = 0;
        pixel_data[125][185] = 0;
        pixel_data[125][186] = 0;
        pixel_data[125][187] = 0;
        pixel_data[125][188] = 0;
        pixel_data[125][189] = 0;
        pixel_data[125][190] = 0;
        pixel_data[125][191] = 0;
        pixel_data[125][192] = 0;
        pixel_data[125][193] = 0;
        pixel_data[125][194] = 0;
        pixel_data[125][195] = 0;
        pixel_data[125][196] = 0;
        pixel_data[125][197] = 0;
        pixel_data[125][198] = 0;
        pixel_data[125][199] = 0; // y=125
        pixel_data[126][0] = 0;
        pixel_data[126][1] = 0;
        pixel_data[126][2] = 0;
        pixel_data[126][3] = 0;
        pixel_data[126][4] = 0;
        pixel_data[126][5] = 0;
        pixel_data[126][6] = 0;
        pixel_data[126][7] = 0;
        pixel_data[126][8] = 0;
        pixel_data[126][9] = 0;
        pixel_data[126][10] = 0;
        pixel_data[126][11] = 0;
        pixel_data[126][12] = 0;
        pixel_data[126][13] = 0;
        pixel_data[126][14] = 0;
        pixel_data[126][15] = 0;
        pixel_data[126][16] = 0;
        pixel_data[126][17] = 0;
        pixel_data[126][18] = 0;
        pixel_data[126][19] = 0;
        pixel_data[126][20] = 0;
        pixel_data[126][21] = 0;
        pixel_data[126][22] = 0;
        pixel_data[126][23] = 0;
        pixel_data[126][24] = 0;
        pixel_data[126][25] = 0;
        pixel_data[126][26] = 0;
        pixel_data[126][27] = 0;
        pixel_data[126][28] = 0;
        pixel_data[126][29] = 0;
        pixel_data[126][30] = 0;
        pixel_data[126][31] = 0;
        pixel_data[126][32] = 0;
        pixel_data[126][33] = 0;
        pixel_data[126][34] = 0;
        pixel_data[126][35] = 0;
        pixel_data[126][36] = 0;
        pixel_data[126][37] = 0;
        pixel_data[126][38] = 0;
        pixel_data[126][39] = 0;
        pixel_data[126][40] = 0;
        pixel_data[126][41] = 0;
        pixel_data[126][42] = 0;
        pixel_data[126][43] = 0;
        pixel_data[126][44] = 0;
        pixel_data[126][45] = 0;
        pixel_data[126][46] = 0;
        pixel_data[126][47] = 0;
        pixel_data[126][48] = 0;
        pixel_data[126][49] = 0;
        pixel_data[126][50] = 0;
        pixel_data[126][51] = 0;
        pixel_data[126][52] = 0;
        pixel_data[126][53] = 0;
        pixel_data[126][54] = 0;
        pixel_data[126][55] = 0;
        pixel_data[126][56] = 0;
        pixel_data[126][57] = 0;
        pixel_data[126][58] = 0;
        pixel_data[126][59] = 0;
        pixel_data[126][60] = 0;
        pixel_data[126][61] = 0;
        pixel_data[126][62] = 0;
        pixel_data[126][63] = 0;
        pixel_data[126][64] = 0;
        pixel_data[126][65] = 0;
        pixel_data[126][66] = 0;
        pixel_data[126][67] = 0;
        pixel_data[126][68] = 0;
        pixel_data[126][69] = 0;
        pixel_data[126][70] = 0;
        pixel_data[126][71] = 0;
        pixel_data[126][72] = 0;
        pixel_data[126][73] = 0;
        pixel_data[126][74] = 0;
        pixel_data[126][75] = 0;
        pixel_data[126][76] = 0;
        pixel_data[126][77] = 0;
        pixel_data[126][78] = 0;
        pixel_data[126][79] = 0;
        pixel_data[126][80] = 0;
        pixel_data[126][81] = 0;
        pixel_data[126][82] = 0;
        pixel_data[126][83] = 0;
        pixel_data[126][84] = 0;
        pixel_data[126][85] = 0;
        pixel_data[126][86] = 0;
        pixel_data[126][87] = 0;
        pixel_data[126][88] = 0;
        pixel_data[126][89] = 0;
        pixel_data[126][90] = 0;
        pixel_data[126][91] = 0;
        pixel_data[126][92] = 0;
        pixel_data[126][93] = 0;
        pixel_data[126][94] = 0;
        pixel_data[126][95] = 0;
        pixel_data[126][96] = 0;
        pixel_data[126][97] = 0;
        pixel_data[126][98] = 0;
        pixel_data[126][99] = 0;
        pixel_data[126][100] = 0;
        pixel_data[126][101] = 0;
        pixel_data[126][102] = 0;
        pixel_data[126][103] = 0;
        pixel_data[126][104] = 0;
        pixel_data[126][105] = 0;
        pixel_data[126][106] = 0;
        pixel_data[126][107] = 0;
        pixel_data[126][108] = 0;
        pixel_data[126][109] = 0;
        pixel_data[126][110] = 0;
        pixel_data[126][111] = 0;
        pixel_data[126][112] = 0;
        pixel_data[126][113] = 0;
        pixel_data[126][114] = 0;
        pixel_data[126][115] = 0;
        pixel_data[126][116] = 0;
        pixel_data[126][117] = 0;
        pixel_data[126][118] = 0;
        pixel_data[126][119] = 0;
        pixel_data[126][120] = 0;
        pixel_data[126][121] = 0;
        pixel_data[126][122] = 0;
        pixel_data[126][123] = 0;
        pixel_data[126][124] = 0;
        pixel_data[126][125] = 0;
        pixel_data[126][126] = 0;
        pixel_data[126][127] = 0;
        pixel_data[126][128] = 0;
        pixel_data[126][129] = 0;
        pixel_data[126][130] = 0;
        pixel_data[126][131] = 0;
        pixel_data[126][132] = 0;
        pixel_data[126][133] = 0;
        pixel_data[126][134] = 0;
        pixel_data[126][135] = 0;
        pixel_data[126][136] = 0;
        pixel_data[126][137] = 0;
        pixel_data[126][138] = 0;
        pixel_data[126][139] = 0;
        pixel_data[126][140] = 0;
        pixel_data[126][141] = 0;
        pixel_data[126][142] = 0;
        pixel_data[126][143] = 0;
        pixel_data[126][144] = 0;
        pixel_data[126][145] = 0;
        pixel_data[126][146] = 0;
        pixel_data[126][147] = 0;
        pixel_data[126][148] = 0;
        pixel_data[126][149] = 0;
        pixel_data[126][150] = 0;
        pixel_data[126][151] = 0;
        pixel_data[126][152] = 0;
        pixel_data[126][153] = 0;
        pixel_data[126][154] = 0;
        pixel_data[126][155] = 0;
        pixel_data[126][156] = 0;
        pixel_data[126][157] = 0;
        pixel_data[126][158] = 0;
        pixel_data[126][159] = 0;
        pixel_data[126][160] = 0;
        pixel_data[126][161] = 0;
        pixel_data[126][162] = 0;
        pixel_data[126][163] = 0;
        pixel_data[126][164] = 0;
        pixel_data[126][165] = 0;
        pixel_data[126][166] = 0;
        pixel_data[126][167] = 0;
        pixel_data[126][168] = 0;
        pixel_data[126][169] = 0;
        pixel_data[126][170] = 0;
        pixel_data[126][171] = 0;
        pixel_data[126][172] = 0;
        pixel_data[126][173] = 0;
        pixel_data[126][174] = 0;
        pixel_data[126][175] = 0;
        pixel_data[126][176] = 0;
        pixel_data[126][177] = 0;
        pixel_data[126][178] = 0;
        pixel_data[126][179] = 0;
        pixel_data[126][180] = 0;
        pixel_data[126][181] = 0;
        pixel_data[126][182] = 0;
        pixel_data[126][183] = 0;
        pixel_data[126][184] = 0;
        pixel_data[126][185] = 0;
        pixel_data[126][186] = 0;
        pixel_data[126][187] = 0;
        pixel_data[126][188] = 0;
        pixel_data[126][189] = 0;
        pixel_data[126][190] = 0;
        pixel_data[126][191] = 0;
        pixel_data[126][192] = 0;
        pixel_data[126][193] = 0;
        pixel_data[126][194] = 0;
        pixel_data[126][195] = 0;
        pixel_data[126][196] = 0;
        pixel_data[126][197] = 0;
        pixel_data[126][198] = 0;
        pixel_data[126][199] = 0; // y=126
        pixel_data[127][0] = 0;
        pixel_data[127][1] = 0;
        pixel_data[127][2] = 0;
        pixel_data[127][3] = 0;
        pixel_data[127][4] = 0;
        pixel_data[127][5] = 0;
        pixel_data[127][6] = 0;
        pixel_data[127][7] = 0;
        pixel_data[127][8] = 0;
        pixel_data[127][9] = 0;
        pixel_data[127][10] = 0;
        pixel_data[127][11] = 0;
        pixel_data[127][12] = 0;
        pixel_data[127][13] = 0;
        pixel_data[127][14] = 0;
        pixel_data[127][15] = 0;
        pixel_data[127][16] = 0;
        pixel_data[127][17] = 0;
        pixel_data[127][18] = 0;
        pixel_data[127][19] = 0;
        pixel_data[127][20] = 0;
        pixel_data[127][21] = 0;
        pixel_data[127][22] = 0;
        pixel_data[127][23] = 0;
        pixel_data[127][24] = 0;
        pixel_data[127][25] = 0;
        pixel_data[127][26] = 0;
        pixel_data[127][27] = 0;
        pixel_data[127][28] = 0;
        pixel_data[127][29] = 0;
        pixel_data[127][30] = 0;
        pixel_data[127][31] = 0;
        pixel_data[127][32] = 0;
        pixel_data[127][33] = 0;
        pixel_data[127][34] = 0;
        pixel_data[127][35] = 0;
        pixel_data[127][36] = 0;
        pixel_data[127][37] = 0;
        pixel_data[127][38] = 0;
        pixel_data[127][39] = 0;
        pixel_data[127][40] = 0;
        pixel_data[127][41] = 0;
        pixel_data[127][42] = 0;
        pixel_data[127][43] = 0;
        pixel_data[127][44] = 0;
        pixel_data[127][45] = 0;
        pixel_data[127][46] = 0;
        pixel_data[127][47] = 0;
        pixel_data[127][48] = 0;
        pixel_data[127][49] = 0;
        pixel_data[127][50] = 0;
        pixel_data[127][51] = 0;
        pixel_data[127][52] = 0;
        pixel_data[127][53] = 0;
        pixel_data[127][54] = 0;
        pixel_data[127][55] = 0;
        pixel_data[127][56] = 0;
        pixel_data[127][57] = 0;
        pixel_data[127][58] = 0;
        pixel_data[127][59] = 0;
        pixel_data[127][60] = 0;
        pixel_data[127][61] = 0;
        pixel_data[127][62] = 0;
        pixel_data[127][63] = 0;
        pixel_data[127][64] = 0;
        pixel_data[127][65] = 0;
        pixel_data[127][66] = 0;
        pixel_data[127][67] = 0;
        pixel_data[127][68] = 0;
        pixel_data[127][69] = 0;
        pixel_data[127][70] = 0;
        pixel_data[127][71] = 0;
        pixel_data[127][72] = 0;
        pixel_data[127][73] = 0;
        pixel_data[127][74] = 0;
        pixel_data[127][75] = 0;
        pixel_data[127][76] = 0;
        pixel_data[127][77] = 0;
        pixel_data[127][78] = 0;
        pixel_data[127][79] = 0;
        pixel_data[127][80] = 0;
        pixel_data[127][81] = 0;
        pixel_data[127][82] = 0;
        pixel_data[127][83] = 0;
        pixel_data[127][84] = 0;
        pixel_data[127][85] = 0;
        pixel_data[127][86] = 0;
        pixel_data[127][87] = 0;
        pixel_data[127][88] = 0;
        pixel_data[127][89] = 0;
        pixel_data[127][90] = 0;
        pixel_data[127][91] = 0;
        pixel_data[127][92] = 0;
        pixel_data[127][93] = 0;
        pixel_data[127][94] = 0;
        pixel_data[127][95] = 0;
        pixel_data[127][96] = 0;
        pixel_data[127][97] = 0;
        pixel_data[127][98] = 0;
        pixel_data[127][99] = 0;
        pixel_data[127][100] = 0;
        pixel_data[127][101] = 0;
        pixel_data[127][102] = 0;
        pixel_data[127][103] = 0;
        pixel_data[127][104] = 0;
        pixel_data[127][105] = 0;
        pixel_data[127][106] = 0;
        pixel_data[127][107] = 0;
        pixel_data[127][108] = 0;
        pixel_data[127][109] = 0;
        pixel_data[127][110] = 0;
        pixel_data[127][111] = 0;
        pixel_data[127][112] = 0;
        pixel_data[127][113] = 0;
        pixel_data[127][114] = 0;
        pixel_data[127][115] = 0;
        pixel_data[127][116] = 0;
        pixel_data[127][117] = 0;
        pixel_data[127][118] = 0;
        pixel_data[127][119] = 0;
        pixel_data[127][120] = 0;
        pixel_data[127][121] = 0;
        pixel_data[127][122] = 0;
        pixel_data[127][123] = 0;
        pixel_data[127][124] = 0;
        pixel_data[127][125] = 0;
        pixel_data[127][126] = 0;
        pixel_data[127][127] = 0;
        pixel_data[127][128] = 0;
        pixel_data[127][129] = 0;
        pixel_data[127][130] = 0;
        pixel_data[127][131] = 0;
        pixel_data[127][132] = 0;
        pixel_data[127][133] = 0;
        pixel_data[127][134] = 0;
        pixel_data[127][135] = 0;
        pixel_data[127][136] = 0;
        pixel_data[127][137] = 0;
        pixel_data[127][138] = 0;
        pixel_data[127][139] = 0;
        pixel_data[127][140] = 0;
        pixel_data[127][141] = 0;
        pixel_data[127][142] = 0;
        pixel_data[127][143] = 0;
        pixel_data[127][144] = 0;
        pixel_data[127][145] = 0;
        pixel_data[127][146] = 0;
        pixel_data[127][147] = 0;
        pixel_data[127][148] = 0;
        pixel_data[127][149] = 0;
        pixel_data[127][150] = 0;
        pixel_data[127][151] = 0;
        pixel_data[127][152] = 0;
        pixel_data[127][153] = 0;
        pixel_data[127][154] = 0;
        pixel_data[127][155] = 0;
        pixel_data[127][156] = 0;
        pixel_data[127][157] = 0;
        pixel_data[127][158] = 0;
        pixel_data[127][159] = 0;
        pixel_data[127][160] = 0;
        pixel_data[127][161] = 0;
        pixel_data[127][162] = 0;
        pixel_data[127][163] = 0;
        pixel_data[127][164] = 0;
        pixel_data[127][165] = 0;
        pixel_data[127][166] = 0;
        pixel_data[127][167] = 0;
        pixel_data[127][168] = 0;
        pixel_data[127][169] = 0;
        pixel_data[127][170] = 0;
        pixel_data[127][171] = 0;
        pixel_data[127][172] = 0;
        pixel_data[127][173] = 0;
        pixel_data[127][174] = 0;
        pixel_data[127][175] = 0;
        pixel_data[127][176] = 0;
        pixel_data[127][177] = 0;
        pixel_data[127][178] = 0;
        pixel_data[127][179] = 0;
        pixel_data[127][180] = 0;
        pixel_data[127][181] = 0;
        pixel_data[127][182] = 0;
        pixel_data[127][183] = 0;
        pixel_data[127][184] = 0;
        pixel_data[127][185] = 0;
        pixel_data[127][186] = 0;
        pixel_data[127][187] = 0;
        pixel_data[127][188] = 0;
        pixel_data[127][189] = 0;
        pixel_data[127][190] = 0;
        pixel_data[127][191] = 0;
        pixel_data[127][192] = 0;
        pixel_data[127][193] = 0;
        pixel_data[127][194] = 0;
        pixel_data[127][195] = 0;
        pixel_data[127][196] = 0;
        pixel_data[127][197] = 0;
        pixel_data[127][198] = 0;
        pixel_data[127][199] = 0; // y=127
        pixel_data[128][0] = 0;
        pixel_data[128][1] = 0;
        pixel_data[128][2] = 0;
        pixel_data[128][3] = 0;
        pixel_data[128][4] = 0;
        pixel_data[128][5] = 0;
        pixel_data[128][6] = 0;
        pixel_data[128][7] = 0;
        pixel_data[128][8] = 0;
        pixel_data[128][9] = 0;
        pixel_data[128][10] = 0;
        pixel_data[128][11] = 0;
        pixel_data[128][12] = 0;
        pixel_data[128][13] = 0;
        pixel_data[128][14] = 0;
        pixel_data[128][15] = 0;
        pixel_data[128][16] = 0;
        pixel_data[128][17] = 0;
        pixel_data[128][18] = 0;
        pixel_data[128][19] = 0;
        pixel_data[128][20] = 0;
        pixel_data[128][21] = 0;
        pixel_data[128][22] = 0;
        pixel_data[128][23] = 0;
        pixel_data[128][24] = 0;
        pixel_data[128][25] = 0;
        pixel_data[128][26] = 0;
        pixel_data[128][27] = 0;
        pixel_data[128][28] = 0;
        pixel_data[128][29] = 0;
        pixel_data[128][30] = 0;
        pixel_data[128][31] = 0;
        pixel_data[128][32] = 0;
        pixel_data[128][33] = 0;
        pixel_data[128][34] = 0;
        pixel_data[128][35] = 0;
        pixel_data[128][36] = 0;
        pixel_data[128][37] = 0;
        pixel_data[128][38] = 0;
        pixel_data[128][39] = 0;
        pixel_data[128][40] = 0;
        pixel_data[128][41] = 0;
        pixel_data[128][42] = 0;
        pixel_data[128][43] = 0;
        pixel_data[128][44] = 0;
        pixel_data[128][45] = 0;
        pixel_data[128][46] = 0;
        pixel_data[128][47] = 0;
        pixel_data[128][48] = 0;
        pixel_data[128][49] = 0;
        pixel_data[128][50] = 0;
        pixel_data[128][51] = 0;
        pixel_data[128][52] = 0;
        pixel_data[128][53] = 0;
        pixel_data[128][54] = 0;
        pixel_data[128][55] = 0;
        pixel_data[128][56] = 0;
        pixel_data[128][57] = 0;
        pixel_data[128][58] = 0;
        pixel_data[128][59] = 0;
        pixel_data[128][60] = 0;
        pixel_data[128][61] = 0;
        pixel_data[128][62] = 0;
        pixel_data[128][63] = 0;
        pixel_data[128][64] = 0;
        pixel_data[128][65] = 0;
        pixel_data[128][66] = 0;
        pixel_data[128][67] = 0;
        pixel_data[128][68] = 0;
        pixel_data[128][69] = 0;
        pixel_data[128][70] = 0;
        pixel_data[128][71] = 0;
        pixel_data[128][72] = 0;
        pixel_data[128][73] = 0;
        pixel_data[128][74] = 0;
        pixel_data[128][75] = 0;
        pixel_data[128][76] = 0;
        pixel_data[128][77] = 0;
        pixel_data[128][78] = 0;
        pixel_data[128][79] = 0;
        pixel_data[128][80] = 0;
        pixel_data[128][81] = 0;
        pixel_data[128][82] = 0;
        pixel_data[128][83] = 0;
        pixel_data[128][84] = 0;
        pixel_data[128][85] = 0;
        pixel_data[128][86] = 0;
        pixel_data[128][87] = 0;
        pixel_data[128][88] = 0;
        pixel_data[128][89] = 0;
        pixel_data[128][90] = 0;
        pixel_data[128][91] = 0;
        pixel_data[128][92] = 0;
        pixel_data[128][93] = 0;
        pixel_data[128][94] = 0;
        pixel_data[128][95] = 0;
        pixel_data[128][96] = 0;
        pixel_data[128][97] = 0;
        pixel_data[128][98] = 0;
        pixel_data[128][99] = 0;
        pixel_data[128][100] = 0;
        pixel_data[128][101] = 0;
        pixel_data[128][102] = 0;
        pixel_data[128][103] = 0;
        pixel_data[128][104] = 0;
        pixel_data[128][105] = 0;
        pixel_data[128][106] = 0;
        pixel_data[128][107] = 0;
        pixel_data[128][108] = 0;
        pixel_data[128][109] = 0;
        pixel_data[128][110] = 0;
        pixel_data[128][111] = 0;
        pixel_data[128][112] = 0;
        pixel_data[128][113] = 0;
        pixel_data[128][114] = 0;
        pixel_data[128][115] = 0;
        pixel_data[128][116] = 0;
        pixel_data[128][117] = 0;
        pixel_data[128][118] = 0;
        pixel_data[128][119] = 0;
        pixel_data[128][120] = 0;
        pixel_data[128][121] = 0;
        pixel_data[128][122] = 0;
        pixel_data[128][123] = 0;
        pixel_data[128][124] = 0;
        pixel_data[128][125] = 0;
        pixel_data[128][126] = 0;
        pixel_data[128][127] = 0;
        pixel_data[128][128] = 0;
        pixel_data[128][129] = 0;
        pixel_data[128][130] = 0;
        pixel_data[128][131] = 0;
        pixel_data[128][132] = 0;
        pixel_data[128][133] = 0;
        pixel_data[128][134] = 0;
        pixel_data[128][135] = 0;
        pixel_data[128][136] = 0;
        pixel_data[128][137] = 0;
        pixel_data[128][138] = 0;
        pixel_data[128][139] = 0;
        pixel_data[128][140] = 0;
        pixel_data[128][141] = 0;
        pixel_data[128][142] = 0;
        pixel_data[128][143] = 0;
        pixel_data[128][144] = 0;
        pixel_data[128][145] = 0;
        pixel_data[128][146] = 0;
        pixel_data[128][147] = 0;
        pixel_data[128][148] = 0;
        pixel_data[128][149] = 0;
        pixel_data[128][150] = 0;
        pixel_data[128][151] = 0;
        pixel_data[128][152] = 0;
        pixel_data[128][153] = 0;
        pixel_data[128][154] = 0;
        pixel_data[128][155] = 0;
        pixel_data[128][156] = 0;
        pixel_data[128][157] = 0;
        pixel_data[128][158] = 0;
        pixel_data[128][159] = 0;
        pixel_data[128][160] = 0;
        pixel_data[128][161] = 0;
        pixel_data[128][162] = 0;
        pixel_data[128][163] = 0;
        pixel_data[128][164] = 0;
        pixel_data[128][165] = 0;
        pixel_data[128][166] = 0;
        pixel_data[128][167] = 0;
        pixel_data[128][168] = 0;
        pixel_data[128][169] = 0;
        pixel_data[128][170] = 0;
        pixel_data[128][171] = 0;
        pixel_data[128][172] = 0;
        pixel_data[128][173] = 0;
        pixel_data[128][174] = 0;
        pixel_data[128][175] = 0;
        pixel_data[128][176] = 0;
        pixel_data[128][177] = 0;
        pixel_data[128][178] = 0;
        pixel_data[128][179] = 0;
        pixel_data[128][180] = 0;
        pixel_data[128][181] = 0;
        pixel_data[128][182] = 0;
        pixel_data[128][183] = 0;
        pixel_data[128][184] = 0;
        pixel_data[128][185] = 0;
        pixel_data[128][186] = 0;
        pixel_data[128][187] = 0;
        pixel_data[128][188] = 0;
        pixel_data[128][189] = 0;
        pixel_data[128][190] = 0;
        pixel_data[128][191] = 0;
        pixel_data[128][192] = 0;
        pixel_data[128][193] = 0;
        pixel_data[128][194] = 0;
        pixel_data[128][195] = 0;
        pixel_data[128][196] = 0;
        pixel_data[128][197] = 0;
        pixel_data[128][198] = 0;
        pixel_data[128][199] = 0; // y=128
        pixel_data[129][0] = 0;
        pixel_data[129][1] = 0;
        pixel_data[129][2] = 0;
        pixel_data[129][3] = 0;
        pixel_data[129][4] = 0;
        pixel_data[129][5] = 0;
        pixel_data[129][6] = 0;
        pixel_data[129][7] = 0;
        pixel_data[129][8] = 0;
        pixel_data[129][9] = 0;
        pixel_data[129][10] = 0;
        pixel_data[129][11] = 0;
        pixel_data[129][12] = 0;
        pixel_data[129][13] = 0;
        pixel_data[129][14] = 0;
        pixel_data[129][15] = 0;
        pixel_data[129][16] = 0;
        pixel_data[129][17] = 0;
        pixel_data[129][18] = 0;
        pixel_data[129][19] = 0;
        pixel_data[129][20] = 0;
        pixel_data[129][21] = 0;
        pixel_data[129][22] = 0;
        pixel_data[129][23] = 0;
        pixel_data[129][24] = 0;
        pixel_data[129][25] = 0;
        pixel_data[129][26] = 0;
        pixel_data[129][27] = 0;
        pixel_data[129][28] = 0;
        pixel_data[129][29] = 0;
        pixel_data[129][30] = 0;
        pixel_data[129][31] = 0;
        pixel_data[129][32] = 0;
        pixel_data[129][33] = 0;
        pixel_data[129][34] = 0;
        pixel_data[129][35] = 0;
        pixel_data[129][36] = 0;
        pixel_data[129][37] = 0;
        pixel_data[129][38] = 0;
        pixel_data[129][39] = 0;
        pixel_data[129][40] = 0;
        pixel_data[129][41] = 0;
        pixel_data[129][42] = 0;
        pixel_data[129][43] = 0;
        pixel_data[129][44] = 0;
        pixel_data[129][45] = 0;
        pixel_data[129][46] = 0;
        pixel_data[129][47] = 0;
        pixel_data[129][48] = 0;
        pixel_data[129][49] = 0;
        pixel_data[129][50] = 0;
        pixel_data[129][51] = 0;
        pixel_data[129][52] = 0;
        pixel_data[129][53] = 0;
        pixel_data[129][54] = 0;
        pixel_data[129][55] = 0;
        pixel_data[129][56] = 0;
        pixel_data[129][57] = 0;
        pixel_data[129][58] = 0;
        pixel_data[129][59] = 0;
        pixel_data[129][60] = 0;
        pixel_data[129][61] = 0;
        pixel_data[129][62] = 0;
        pixel_data[129][63] = 0;
        pixel_data[129][64] = 0;
        pixel_data[129][65] = 0;
        pixel_data[129][66] = 0;
        pixel_data[129][67] = 0;
        pixel_data[129][68] = 0;
        pixel_data[129][69] = 0;
        pixel_data[129][70] = 0;
        pixel_data[129][71] = 0;
        pixel_data[129][72] = 0;
        pixel_data[129][73] = 0;
        pixel_data[129][74] = 0;
        pixel_data[129][75] = 0;
        pixel_data[129][76] = 0;
        pixel_data[129][77] = 0;
        pixel_data[129][78] = 0;
        pixel_data[129][79] = 0;
        pixel_data[129][80] = 0;
        pixel_data[129][81] = 0;
        pixel_data[129][82] = 0;
        pixel_data[129][83] = 0;
        pixel_data[129][84] = 0;
        pixel_data[129][85] = 0;
        pixel_data[129][86] = 0;
        pixel_data[129][87] = 0;
        pixel_data[129][88] = 0;
        pixel_data[129][89] = 0;
        pixel_data[129][90] = 0;
        pixel_data[129][91] = 0;
        pixel_data[129][92] = 0;
        pixel_data[129][93] = 0;
        pixel_data[129][94] = 0;
        pixel_data[129][95] = 0;
        pixel_data[129][96] = 0;
        pixel_data[129][97] = 0;
        pixel_data[129][98] = 0;
        pixel_data[129][99] = 0;
        pixel_data[129][100] = 0;
        pixel_data[129][101] = 0;
        pixel_data[129][102] = 0;
        pixel_data[129][103] = 0;
        pixel_data[129][104] = 0;
        pixel_data[129][105] = 0;
        pixel_data[129][106] = 0;
        pixel_data[129][107] = 0;
        pixel_data[129][108] = 0;
        pixel_data[129][109] = 0;
        pixel_data[129][110] = 0;
        pixel_data[129][111] = 0;
        pixel_data[129][112] = 0;
        pixel_data[129][113] = 0;
        pixel_data[129][114] = 0;
        pixel_data[129][115] = 0;
        pixel_data[129][116] = 0;
        pixel_data[129][117] = 0;
        pixel_data[129][118] = 0;
        pixel_data[129][119] = 0;
        pixel_data[129][120] = 0;
        pixel_data[129][121] = 0;
        pixel_data[129][122] = 0;
        pixel_data[129][123] = 0;
        pixel_data[129][124] = 0;
        pixel_data[129][125] = 0;
        pixel_data[129][126] = 0;
        pixel_data[129][127] = 0;
        pixel_data[129][128] = 0;
        pixel_data[129][129] = 0;
        pixel_data[129][130] = 0;
        pixel_data[129][131] = 0;
        pixel_data[129][132] = 0;
        pixel_data[129][133] = 0;
        pixel_data[129][134] = 0;
        pixel_data[129][135] = 0;
        pixel_data[129][136] = 0;
        pixel_data[129][137] = 0;
        pixel_data[129][138] = 0;
        pixel_data[129][139] = 0;
        pixel_data[129][140] = 0;
        pixel_data[129][141] = 0;
        pixel_data[129][142] = 0;
        pixel_data[129][143] = 0;
        pixel_data[129][144] = 0;
        pixel_data[129][145] = 0;
        pixel_data[129][146] = 0;
        pixel_data[129][147] = 0;
        pixel_data[129][148] = 0;
        pixel_data[129][149] = 0;
        pixel_data[129][150] = 0;
        pixel_data[129][151] = 0;
        pixel_data[129][152] = 0;
        pixel_data[129][153] = 0;
        pixel_data[129][154] = 0;
        pixel_data[129][155] = 0;
        pixel_data[129][156] = 0;
        pixel_data[129][157] = 0;
        pixel_data[129][158] = 0;
        pixel_data[129][159] = 0;
        pixel_data[129][160] = 0;
        pixel_data[129][161] = 0;
        pixel_data[129][162] = 0;
        pixel_data[129][163] = 0;
        pixel_data[129][164] = 0;
        pixel_data[129][165] = 0;
        pixel_data[129][166] = 0;
        pixel_data[129][167] = 0;
        pixel_data[129][168] = 0;
        pixel_data[129][169] = 0;
        pixel_data[129][170] = 0;
        pixel_data[129][171] = 0;
        pixel_data[129][172] = 0;
        pixel_data[129][173] = 0;
        pixel_data[129][174] = 0;
        pixel_data[129][175] = 0;
        pixel_data[129][176] = 0;
        pixel_data[129][177] = 0;
        pixel_data[129][178] = 0;
        pixel_data[129][179] = 0;
        pixel_data[129][180] = 0;
        pixel_data[129][181] = 0;
        pixel_data[129][182] = 0;
        pixel_data[129][183] = 0;
        pixel_data[129][184] = 0;
        pixel_data[129][185] = 0;
        pixel_data[129][186] = 0;
        pixel_data[129][187] = 0;
        pixel_data[129][188] = 0;
        pixel_data[129][189] = 0;
        pixel_data[129][190] = 0;
        pixel_data[129][191] = 0;
        pixel_data[129][192] = 0;
        pixel_data[129][193] = 0;
        pixel_data[129][194] = 0;
        pixel_data[129][195] = 0;
        pixel_data[129][196] = 0;
        pixel_data[129][197] = 0;
        pixel_data[129][198] = 0;
        pixel_data[129][199] = 0; // y=129
        pixel_data[130][0] = 0;
        pixel_data[130][1] = 0;
        pixel_data[130][2] = 0;
        pixel_data[130][3] = 0;
        pixel_data[130][4] = 0;
        pixel_data[130][5] = 0;
        pixel_data[130][6] = 0;
        pixel_data[130][7] = 0;
        pixel_data[130][8] = 0;
        pixel_data[130][9] = 0;
        pixel_data[130][10] = 0;
        pixel_data[130][11] = 0;
        pixel_data[130][12] = 0;
        pixel_data[130][13] = 0;
        pixel_data[130][14] = 0;
        pixel_data[130][15] = 0;
        pixel_data[130][16] = 0;
        pixel_data[130][17] = 0;
        pixel_data[130][18] = 0;
        pixel_data[130][19] = 0;
        pixel_data[130][20] = 0;
        pixel_data[130][21] = 0;
        pixel_data[130][22] = 0;
        pixel_data[130][23] = 0;
        pixel_data[130][24] = 0;
        pixel_data[130][25] = 0;
        pixel_data[130][26] = 0;
        pixel_data[130][27] = 0;
        pixel_data[130][28] = 0;
        pixel_data[130][29] = 0;
        pixel_data[130][30] = 0;
        pixel_data[130][31] = 0;
        pixel_data[130][32] = 0;
        pixel_data[130][33] = 0;
        pixel_data[130][34] = 0;
        pixel_data[130][35] = 0;
        pixel_data[130][36] = 0;
        pixel_data[130][37] = 0;
        pixel_data[130][38] = 0;
        pixel_data[130][39] = 0;
        pixel_data[130][40] = 0;
        pixel_data[130][41] = 0;
        pixel_data[130][42] = 0;
        pixel_data[130][43] = 0;
        pixel_data[130][44] = 0;
        pixel_data[130][45] = 0;
        pixel_data[130][46] = 0;
        pixel_data[130][47] = 0;
        pixel_data[130][48] = 0;
        pixel_data[130][49] = 0;
        pixel_data[130][50] = 0;
        pixel_data[130][51] = 0;
        pixel_data[130][52] = 0;
        pixel_data[130][53] = 0;
        pixel_data[130][54] = 0;
        pixel_data[130][55] = 0;
        pixel_data[130][56] = 0;
        pixel_data[130][57] = 0;
        pixel_data[130][58] = 0;
        pixel_data[130][59] = 0;
        pixel_data[130][60] = 0;
        pixel_data[130][61] = 0;
        pixel_data[130][62] = 0;
        pixel_data[130][63] = 0;
        pixel_data[130][64] = 0;
        pixel_data[130][65] = 0;
        pixel_data[130][66] = 0;
        pixel_data[130][67] = 0;
        pixel_data[130][68] = 0;
        pixel_data[130][69] = 0;
        pixel_data[130][70] = 0;
        pixel_data[130][71] = 0;
        pixel_data[130][72] = 0;
        pixel_data[130][73] = 0;
        pixel_data[130][74] = 0;
        pixel_data[130][75] = 0;
        pixel_data[130][76] = 0;
        pixel_data[130][77] = 0;
        pixel_data[130][78] = 0;
        pixel_data[130][79] = 0;
        pixel_data[130][80] = 0;
        pixel_data[130][81] = 0;
        pixel_data[130][82] = 0;
        pixel_data[130][83] = 0;
        pixel_data[130][84] = 0;
        pixel_data[130][85] = 0;
        pixel_data[130][86] = 0;
        pixel_data[130][87] = 0;
        pixel_data[130][88] = 0;
        pixel_data[130][89] = 0;
        pixel_data[130][90] = 0;
        pixel_data[130][91] = 0;
        pixel_data[130][92] = 0;
        pixel_data[130][93] = 0;
        pixel_data[130][94] = 0;
        pixel_data[130][95] = 0;
        pixel_data[130][96] = 0;
        pixel_data[130][97] = 0;
        pixel_data[130][98] = 0;
        pixel_data[130][99] = 0;
        pixel_data[130][100] = 0;
        pixel_data[130][101] = 0;
        pixel_data[130][102] = 0;
        pixel_data[130][103] = 0;
        pixel_data[130][104] = 0;
        pixel_data[130][105] = 0;
        pixel_data[130][106] = 0;
        pixel_data[130][107] = 0;
        pixel_data[130][108] = 0;
        pixel_data[130][109] = 0;
        pixel_data[130][110] = 0;
        pixel_data[130][111] = 0;
        pixel_data[130][112] = 0;
        pixel_data[130][113] = 0;
        pixel_data[130][114] = 0;
        pixel_data[130][115] = 0;
        pixel_data[130][116] = 0;
        pixel_data[130][117] = 0;
        pixel_data[130][118] = 0;
        pixel_data[130][119] = 0;
        pixel_data[130][120] = 0;
        pixel_data[130][121] = 0;
        pixel_data[130][122] = 0;
        pixel_data[130][123] = 0;
        pixel_data[130][124] = 0;
        pixel_data[130][125] = 0;
        pixel_data[130][126] = 0;
        pixel_data[130][127] = 0;
        pixel_data[130][128] = 0;
        pixel_data[130][129] = 0;
        pixel_data[130][130] = 0;
        pixel_data[130][131] = 0;
        pixel_data[130][132] = 0;
        pixel_data[130][133] = 0;
        pixel_data[130][134] = 0;
        pixel_data[130][135] = 0;
        pixel_data[130][136] = 0;
        pixel_data[130][137] = 0;
        pixel_data[130][138] = 0;
        pixel_data[130][139] = 0;
        pixel_data[130][140] = 0;
        pixel_data[130][141] = 0;
        pixel_data[130][142] = 0;
        pixel_data[130][143] = 0;
        pixel_data[130][144] = 0;
        pixel_data[130][145] = 0;
        pixel_data[130][146] = 0;
        pixel_data[130][147] = 0;
        pixel_data[130][148] = 0;
        pixel_data[130][149] = 0;
        pixel_data[130][150] = 0;
        pixel_data[130][151] = 0;
        pixel_data[130][152] = 0;
        pixel_data[130][153] = 0;
        pixel_data[130][154] = 0;
        pixel_data[130][155] = 0;
        pixel_data[130][156] = 0;
        pixel_data[130][157] = 0;
        pixel_data[130][158] = 0;
        pixel_data[130][159] = 0;
        pixel_data[130][160] = 0;
        pixel_data[130][161] = 0;
        pixel_data[130][162] = 0;
        pixel_data[130][163] = 0;
        pixel_data[130][164] = 0;
        pixel_data[130][165] = 0;
        pixel_data[130][166] = 0;
        pixel_data[130][167] = 0;
        pixel_data[130][168] = 0;
        pixel_data[130][169] = 0;
        pixel_data[130][170] = 0;
        pixel_data[130][171] = 0;
        pixel_data[130][172] = 0;
        pixel_data[130][173] = 0;
        pixel_data[130][174] = 0;
        pixel_data[130][175] = 0;
        pixel_data[130][176] = 0;
        pixel_data[130][177] = 0;
        pixel_data[130][178] = 0;
        pixel_data[130][179] = 0;
        pixel_data[130][180] = 0;
        pixel_data[130][181] = 0;
        pixel_data[130][182] = 0;
        pixel_data[130][183] = 0;
        pixel_data[130][184] = 0;
        pixel_data[130][185] = 0;
        pixel_data[130][186] = 0;
        pixel_data[130][187] = 0;
        pixel_data[130][188] = 0;
        pixel_data[130][189] = 0;
        pixel_data[130][190] = 0;
        pixel_data[130][191] = 0;
        pixel_data[130][192] = 0;
        pixel_data[130][193] = 0;
        pixel_data[130][194] = 0;
        pixel_data[130][195] = 0;
        pixel_data[130][196] = 0;
        pixel_data[130][197] = 0;
        pixel_data[130][198] = 0;
        pixel_data[130][199] = 0; // y=130
        pixel_data[131][0] = 0;
        pixel_data[131][1] = 0;
        pixel_data[131][2] = 0;
        pixel_data[131][3] = 0;
        pixel_data[131][4] = 0;
        pixel_data[131][5] = 0;
        pixel_data[131][6] = 0;
        pixel_data[131][7] = 0;
        pixel_data[131][8] = 0;
        pixel_data[131][9] = 0;
        pixel_data[131][10] = 0;
        pixel_data[131][11] = 0;
        pixel_data[131][12] = 0;
        pixel_data[131][13] = 0;
        pixel_data[131][14] = 0;
        pixel_data[131][15] = 0;
        pixel_data[131][16] = 0;
        pixel_data[131][17] = 0;
        pixel_data[131][18] = 0;
        pixel_data[131][19] = 0;
        pixel_data[131][20] = 0;
        pixel_data[131][21] = 0;
        pixel_data[131][22] = 0;
        pixel_data[131][23] = 0;
        pixel_data[131][24] = 0;
        pixel_data[131][25] = 0;
        pixel_data[131][26] = 0;
        pixel_data[131][27] = 0;
        pixel_data[131][28] = 0;
        pixel_data[131][29] = 0;
        pixel_data[131][30] = 0;
        pixel_data[131][31] = 0;
        pixel_data[131][32] = 0;
        pixel_data[131][33] = 0;
        pixel_data[131][34] = 0;
        pixel_data[131][35] = 0;
        pixel_data[131][36] = 0;
        pixel_data[131][37] = 0;
        pixel_data[131][38] = 0;
        pixel_data[131][39] = 0;
        pixel_data[131][40] = 0;
        pixel_data[131][41] = 0;
        pixel_data[131][42] = 0;
        pixel_data[131][43] = 0;
        pixel_data[131][44] = 0;
        pixel_data[131][45] = 0;
        pixel_data[131][46] = 0;
        pixel_data[131][47] = 0;
        pixel_data[131][48] = 0;
        pixel_data[131][49] = 0;
        pixel_data[131][50] = 0;
        pixel_data[131][51] = 0;
        pixel_data[131][52] = 0;
        pixel_data[131][53] = 0;
        pixel_data[131][54] = 0;
        pixel_data[131][55] = 0;
        pixel_data[131][56] = 0;
        pixel_data[131][57] = 0;
        pixel_data[131][58] = 0;
        pixel_data[131][59] = 0;
        pixel_data[131][60] = 0;
        pixel_data[131][61] = 0;
        pixel_data[131][62] = 0;
        pixel_data[131][63] = 0;
        pixel_data[131][64] = 0;
        pixel_data[131][65] = 0;
        pixel_data[131][66] = 0;
        pixel_data[131][67] = 0;
        pixel_data[131][68] = 0;
        pixel_data[131][69] = 0;
        pixel_data[131][70] = 0;
        pixel_data[131][71] = 0;
        pixel_data[131][72] = 0;
        pixel_data[131][73] = 0;
        pixel_data[131][74] = 0;
        pixel_data[131][75] = 0;
        pixel_data[131][76] = 0;
        pixel_data[131][77] = 0;
        pixel_data[131][78] = 0;
        pixel_data[131][79] = 0;
        pixel_data[131][80] = 0;
        pixel_data[131][81] = 0;
        pixel_data[131][82] = 0;
        pixel_data[131][83] = 0;
        pixel_data[131][84] = 0;
        pixel_data[131][85] = 0;
        pixel_data[131][86] = 0;
        pixel_data[131][87] = 0;
        pixel_data[131][88] = 0;
        pixel_data[131][89] = 0;
        pixel_data[131][90] = 0;
        pixel_data[131][91] = 0;
        pixel_data[131][92] = 0;
        pixel_data[131][93] = 0;
        pixel_data[131][94] = 0;
        pixel_data[131][95] = 0;
        pixel_data[131][96] = 0;
        pixel_data[131][97] = 0;
        pixel_data[131][98] = 0;
        pixel_data[131][99] = 0;
        pixel_data[131][100] = 0;
        pixel_data[131][101] = 0;
        pixel_data[131][102] = 0;
        pixel_data[131][103] = 0;
        pixel_data[131][104] = 0;
        pixel_data[131][105] = 0;
        pixel_data[131][106] = 0;
        pixel_data[131][107] = 0;
        pixel_data[131][108] = 0;
        pixel_data[131][109] = 0;
        pixel_data[131][110] = 0;
        pixel_data[131][111] = 0;
        pixel_data[131][112] = 0;
        pixel_data[131][113] = 0;
        pixel_data[131][114] = 0;
        pixel_data[131][115] = 0;
        pixel_data[131][116] = 0;
        pixel_data[131][117] = 0;
        pixel_data[131][118] = 0;
        pixel_data[131][119] = 0;
        pixel_data[131][120] = 0;
        pixel_data[131][121] = 0;
        pixel_data[131][122] = 0;
        pixel_data[131][123] = 0;
        pixel_data[131][124] = 0;
        pixel_data[131][125] = 0;
        pixel_data[131][126] = 0;
        pixel_data[131][127] = 0;
        pixel_data[131][128] = 0;
        pixel_data[131][129] = 0;
        pixel_data[131][130] = 0;
        pixel_data[131][131] = 0;
        pixel_data[131][132] = 0;
        pixel_data[131][133] = 0;
        pixel_data[131][134] = 0;
        pixel_data[131][135] = 0;
        pixel_data[131][136] = 0;
        pixel_data[131][137] = 0;
        pixel_data[131][138] = 0;
        pixel_data[131][139] = 0;
        pixel_data[131][140] = 0;
        pixel_data[131][141] = 0;
        pixel_data[131][142] = 0;
        pixel_data[131][143] = 0;
        pixel_data[131][144] = 0;
        pixel_data[131][145] = 0;
        pixel_data[131][146] = 0;
        pixel_data[131][147] = 0;
        pixel_data[131][148] = 0;
        pixel_data[131][149] = 0;
        pixel_data[131][150] = 0;
        pixel_data[131][151] = 0;
        pixel_data[131][152] = 0;
        pixel_data[131][153] = 0;
        pixel_data[131][154] = 0;
        pixel_data[131][155] = 0;
        pixel_data[131][156] = 0;
        pixel_data[131][157] = 0;
        pixel_data[131][158] = 0;
        pixel_data[131][159] = 0;
        pixel_data[131][160] = 0;
        pixel_data[131][161] = 0;
        pixel_data[131][162] = 0;
        pixel_data[131][163] = 0;
        pixel_data[131][164] = 0;
        pixel_data[131][165] = 0;
        pixel_data[131][166] = 0;
        pixel_data[131][167] = 0;
        pixel_data[131][168] = 0;
        pixel_data[131][169] = 0;
        pixel_data[131][170] = 0;
        pixel_data[131][171] = 0;
        pixel_data[131][172] = 0;
        pixel_data[131][173] = 0;
        pixel_data[131][174] = 0;
        pixel_data[131][175] = 0;
        pixel_data[131][176] = 0;
        pixel_data[131][177] = 0;
        pixel_data[131][178] = 0;
        pixel_data[131][179] = 0;
        pixel_data[131][180] = 0;
        pixel_data[131][181] = 0;
        pixel_data[131][182] = 0;
        pixel_data[131][183] = 0;
        pixel_data[131][184] = 0;
        pixel_data[131][185] = 0;
        pixel_data[131][186] = 0;
        pixel_data[131][187] = 0;
        pixel_data[131][188] = 0;
        pixel_data[131][189] = 0;
        pixel_data[131][190] = 0;
        pixel_data[131][191] = 0;
        pixel_data[131][192] = 0;
        pixel_data[131][193] = 0;
        pixel_data[131][194] = 0;
        pixel_data[131][195] = 0;
        pixel_data[131][196] = 0;
        pixel_data[131][197] = 0;
        pixel_data[131][198] = 0;
        pixel_data[131][199] = 0; // y=131
        pixel_data[132][0] = 0;
        pixel_data[132][1] = 0;
        pixel_data[132][2] = 0;
        pixel_data[132][3] = 0;
        pixel_data[132][4] = 0;
        pixel_data[132][5] = 0;
        pixel_data[132][6] = 0;
        pixel_data[132][7] = 0;
        pixel_data[132][8] = 0;
        pixel_data[132][9] = 0;
        pixel_data[132][10] = 0;
        pixel_data[132][11] = 0;
        pixel_data[132][12] = 0;
        pixel_data[132][13] = 0;
        pixel_data[132][14] = 0;
        pixel_data[132][15] = 0;
        pixel_data[132][16] = 0;
        pixel_data[132][17] = 0;
        pixel_data[132][18] = 0;
        pixel_data[132][19] = 0;
        pixel_data[132][20] = 0;
        pixel_data[132][21] = 0;
        pixel_data[132][22] = 0;
        pixel_data[132][23] = 0;
        pixel_data[132][24] = 0;
        pixel_data[132][25] = 0;
        pixel_data[132][26] = 0;
        pixel_data[132][27] = 0;
        pixel_data[132][28] = 0;
        pixel_data[132][29] = 0;
        pixel_data[132][30] = 0;
        pixel_data[132][31] = 0;
        pixel_data[132][32] = 0;
        pixel_data[132][33] = 0;
        pixel_data[132][34] = 0;
        pixel_data[132][35] = 0;
        pixel_data[132][36] = 0;
        pixel_data[132][37] = 0;
        pixel_data[132][38] = 0;
        pixel_data[132][39] = 0;
        pixel_data[132][40] = 0;
        pixel_data[132][41] = 0;
        pixel_data[132][42] = 0;
        pixel_data[132][43] = 0;
        pixel_data[132][44] = 0;
        pixel_data[132][45] = 0;
        pixel_data[132][46] = 0;
        pixel_data[132][47] = 0;
        pixel_data[132][48] = 0;
        pixel_data[132][49] = 0;
        pixel_data[132][50] = 0;
        pixel_data[132][51] = 0;
        pixel_data[132][52] = 0;
        pixel_data[132][53] = 0;
        pixel_data[132][54] = 0;
        pixel_data[132][55] = 0;
        pixel_data[132][56] = 0;
        pixel_data[132][57] = 0;
        pixel_data[132][58] = 0;
        pixel_data[132][59] = 0;
        pixel_data[132][60] = 0;
        pixel_data[132][61] = 0;
        pixel_data[132][62] = 0;
        pixel_data[132][63] = 0;
        pixel_data[132][64] = 0;
        pixel_data[132][65] = 0;
        pixel_data[132][66] = 0;
        pixel_data[132][67] = 0;
        pixel_data[132][68] = 0;
        pixel_data[132][69] = 0;
        pixel_data[132][70] = 0;
        pixel_data[132][71] = 0;
        pixel_data[132][72] = 0;
        pixel_data[132][73] = 0;
        pixel_data[132][74] = 0;
        pixel_data[132][75] = 0;
        pixel_data[132][76] = 0;
        pixel_data[132][77] = 0;
        pixel_data[132][78] = 0;
        pixel_data[132][79] = 0;
        pixel_data[132][80] = 0;
        pixel_data[132][81] = 0;
        pixel_data[132][82] = 0;
        pixel_data[132][83] = 0;
        pixel_data[132][84] = 0;
        pixel_data[132][85] = 0;
        pixel_data[132][86] = 0;
        pixel_data[132][87] = 0;
        pixel_data[132][88] = 0;
        pixel_data[132][89] = 0;
        pixel_data[132][90] = 0;
        pixel_data[132][91] = 0;
        pixel_data[132][92] = 0;
        pixel_data[132][93] = 0;
        pixel_data[132][94] = 0;
        pixel_data[132][95] = 0;
        pixel_data[132][96] = 0;
        pixel_data[132][97] = 0;
        pixel_data[132][98] = 0;
        pixel_data[132][99] = 0;
        pixel_data[132][100] = 0;
        pixel_data[132][101] = 0;
        pixel_data[132][102] = 0;
        pixel_data[132][103] = 0;
        pixel_data[132][104] = 0;
        pixel_data[132][105] = 0;
        pixel_data[132][106] = 0;
        pixel_data[132][107] = 0;
        pixel_data[132][108] = 0;
        pixel_data[132][109] = 0;
        pixel_data[132][110] = 0;
        pixel_data[132][111] = 0;
        pixel_data[132][112] = 0;
        pixel_data[132][113] = 0;
        pixel_data[132][114] = 0;
        pixel_data[132][115] = 0;
        pixel_data[132][116] = 0;
        pixel_data[132][117] = 0;
        pixel_data[132][118] = 0;
        pixel_data[132][119] = 0;
        pixel_data[132][120] = 0;
        pixel_data[132][121] = 0;
        pixel_data[132][122] = 0;
        pixel_data[132][123] = 0;
        pixel_data[132][124] = 0;
        pixel_data[132][125] = 0;
        pixel_data[132][126] = 0;
        pixel_data[132][127] = 0;
        pixel_data[132][128] = 0;
        pixel_data[132][129] = 0;
        pixel_data[132][130] = 0;
        pixel_data[132][131] = 0;
        pixel_data[132][132] = 0;
        pixel_data[132][133] = 0;
        pixel_data[132][134] = 0;
        pixel_data[132][135] = 0;
        pixel_data[132][136] = 0;
        pixel_data[132][137] = 0;
        pixel_data[132][138] = 0;
        pixel_data[132][139] = 0;
        pixel_data[132][140] = 0;
        pixel_data[132][141] = 0;
        pixel_data[132][142] = 0;
        pixel_data[132][143] = 0;
        pixel_data[132][144] = 0;
        pixel_data[132][145] = 0;
        pixel_data[132][146] = 0;
        pixel_data[132][147] = 0;
        pixel_data[132][148] = 0;
        pixel_data[132][149] = 0;
        pixel_data[132][150] = 0;
        pixel_data[132][151] = 0;
        pixel_data[132][152] = 0;
        pixel_data[132][153] = 0;
        pixel_data[132][154] = 0;
        pixel_data[132][155] = 0;
        pixel_data[132][156] = 0;
        pixel_data[132][157] = 0;
        pixel_data[132][158] = 0;
        pixel_data[132][159] = 0;
        pixel_data[132][160] = 0;
        pixel_data[132][161] = 0;
        pixel_data[132][162] = 0;
        pixel_data[132][163] = 0;
        pixel_data[132][164] = 0;
        pixel_data[132][165] = 0;
        pixel_data[132][166] = 0;
        pixel_data[132][167] = 0;
        pixel_data[132][168] = 0;
        pixel_data[132][169] = 0;
        pixel_data[132][170] = 0;
        pixel_data[132][171] = 0;
        pixel_data[132][172] = 0;
        pixel_data[132][173] = 0;
        pixel_data[132][174] = 0;
        pixel_data[132][175] = 0;
        pixel_data[132][176] = 0;
        pixel_data[132][177] = 0;
        pixel_data[132][178] = 0;
        pixel_data[132][179] = 0;
        pixel_data[132][180] = 0;
        pixel_data[132][181] = 0;
        pixel_data[132][182] = 0;
        pixel_data[132][183] = 0;
        pixel_data[132][184] = 0;
        pixel_data[132][185] = 0;
        pixel_data[132][186] = 0;
        pixel_data[132][187] = 0;
        pixel_data[132][188] = 0;
        pixel_data[132][189] = 0;
        pixel_data[132][190] = 0;
        pixel_data[132][191] = 0;
        pixel_data[132][192] = 0;
        pixel_data[132][193] = 0;
        pixel_data[132][194] = 0;
        pixel_data[132][195] = 0;
        pixel_data[132][196] = 0;
        pixel_data[132][197] = 0;
        pixel_data[132][198] = 0;
        pixel_data[132][199] = 0; // y=132
        pixel_data[133][0] = 0;
        pixel_data[133][1] = 0;
        pixel_data[133][2] = 0;
        pixel_data[133][3] = 0;
        pixel_data[133][4] = 0;
        pixel_data[133][5] = 0;
        pixel_data[133][6] = 0;
        pixel_data[133][7] = 0;
        pixel_data[133][8] = 0;
        pixel_data[133][9] = 0;
        pixel_data[133][10] = 0;
        pixel_data[133][11] = 0;
        pixel_data[133][12] = 0;
        pixel_data[133][13] = 0;
        pixel_data[133][14] = 0;
        pixel_data[133][15] = 0;
        pixel_data[133][16] = 0;
        pixel_data[133][17] = 0;
        pixel_data[133][18] = 0;
        pixel_data[133][19] = 0;
        pixel_data[133][20] = 0;
        pixel_data[133][21] = 0;
        pixel_data[133][22] = 0;
        pixel_data[133][23] = 0;
        pixel_data[133][24] = 0;
        pixel_data[133][25] = 0;
        pixel_data[133][26] = 0;
        pixel_data[133][27] = 0;
        pixel_data[133][28] = 0;
        pixel_data[133][29] = 0;
        pixel_data[133][30] = 0;
        pixel_data[133][31] = 0;
        pixel_data[133][32] = 0;
        pixel_data[133][33] = 0;
        pixel_data[133][34] = 0;
        pixel_data[133][35] = 0;
        pixel_data[133][36] = 0;
        pixel_data[133][37] = 0;
        pixel_data[133][38] = 0;
        pixel_data[133][39] = 0;
        pixel_data[133][40] = 0;
        pixel_data[133][41] = 0;
        pixel_data[133][42] = 0;
        pixel_data[133][43] = 0;
        pixel_data[133][44] = 0;
        pixel_data[133][45] = 0;
        pixel_data[133][46] = 0;
        pixel_data[133][47] = 0;
        pixel_data[133][48] = 0;
        pixel_data[133][49] = 0;
        pixel_data[133][50] = 0;
        pixel_data[133][51] = 0;
        pixel_data[133][52] = 0;
        pixel_data[133][53] = 0;
        pixel_data[133][54] = 0;
        pixel_data[133][55] = 0;
        pixel_data[133][56] = 0;
        pixel_data[133][57] = 0;
        pixel_data[133][58] = 0;
        pixel_data[133][59] = 0;
        pixel_data[133][60] = 0;
        pixel_data[133][61] = 0;
        pixel_data[133][62] = 0;
        pixel_data[133][63] = 0;
        pixel_data[133][64] = 0;
        pixel_data[133][65] = 0;
        pixel_data[133][66] = 0;
        pixel_data[133][67] = 0;
        pixel_data[133][68] = 0;
        pixel_data[133][69] = 0;
        pixel_data[133][70] = 0;
        pixel_data[133][71] = 0;
        pixel_data[133][72] = 0;
        pixel_data[133][73] = 0;
        pixel_data[133][74] = 0;
        pixel_data[133][75] = 0;
        pixel_data[133][76] = 0;
        pixel_data[133][77] = 0;
        pixel_data[133][78] = 0;
        pixel_data[133][79] = 0;
        pixel_data[133][80] = 0;
        pixel_data[133][81] = 0;
        pixel_data[133][82] = 0;
        pixel_data[133][83] = 0;
        pixel_data[133][84] = 0;
        pixel_data[133][85] = 0;
        pixel_data[133][86] = 0;
        pixel_data[133][87] = 0;
        pixel_data[133][88] = 0;
        pixel_data[133][89] = 0;
        pixel_data[133][90] = 0;
        pixel_data[133][91] = 0;
        pixel_data[133][92] = 0;
        pixel_data[133][93] = 0;
        pixel_data[133][94] = 0;
        pixel_data[133][95] = 0;
        pixel_data[133][96] = 0;
        pixel_data[133][97] = 0;
        pixel_data[133][98] = 0;
        pixel_data[133][99] = 0;
        pixel_data[133][100] = 0;
        pixel_data[133][101] = 0;
        pixel_data[133][102] = 0;
        pixel_data[133][103] = 0;
        pixel_data[133][104] = 0;
        pixel_data[133][105] = 0;
        pixel_data[133][106] = 0;
        pixel_data[133][107] = 0;
        pixel_data[133][108] = 0;
        pixel_data[133][109] = 0;
        pixel_data[133][110] = 0;
        pixel_data[133][111] = 0;
        pixel_data[133][112] = 0;
        pixel_data[133][113] = 0;
        pixel_data[133][114] = 0;
        pixel_data[133][115] = 0;
        pixel_data[133][116] = 0;
        pixel_data[133][117] = 0;
        pixel_data[133][118] = 0;
        pixel_data[133][119] = 0;
        pixel_data[133][120] = 0;
        pixel_data[133][121] = 0;
        pixel_data[133][122] = 0;
        pixel_data[133][123] = 0;
        pixel_data[133][124] = 0;
        pixel_data[133][125] = 0;
        pixel_data[133][126] = 0;
        pixel_data[133][127] = 0;
        pixel_data[133][128] = 0;
        pixel_data[133][129] = 0;
        pixel_data[133][130] = 0;
        pixel_data[133][131] = 0;
        pixel_data[133][132] = 0;
        pixel_data[133][133] = 0;
        pixel_data[133][134] = 0;
        pixel_data[133][135] = 0;
        pixel_data[133][136] = 0;
        pixel_data[133][137] = 0;
        pixel_data[133][138] = 0;
        pixel_data[133][139] = 0;
        pixel_data[133][140] = 0;
        pixel_data[133][141] = 0;
        pixel_data[133][142] = 0;
        pixel_data[133][143] = 0;
        pixel_data[133][144] = 0;
        pixel_data[133][145] = 0;
        pixel_data[133][146] = 0;
        pixel_data[133][147] = 0;
        pixel_data[133][148] = 0;
        pixel_data[133][149] = 0;
        pixel_data[133][150] = 0;
        pixel_data[133][151] = 0;
        pixel_data[133][152] = 0;
        pixel_data[133][153] = 0;
        pixel_data[133][154] = 0;
        pixel_data[133][155] = 0;
        pixel_data[133][156] = 0;
        pixel_data[133][157] = 0;
        pixel_data[133][158] = 0;
        pixel_data[133][159] = 0;
        pixel_data[133][160] = 0;
        pixel_data[133][161] = 0;
        pixel_data[133][162] = 0;
        pixel_data[133][163] = 0;
        pixel_data[133][164] = 0;
        pixel_data[133][165] = 0;
        pixel_data[133][166] = 0;
        pixel_data[133][167] = 0;
        pixel_data[133][168] = 0;
        pixel_data[133][169] = 0;
        pixel_data[133][170] = 0;
        pixel_data[133][171] = 0;
        pixel_data[133][172] = 0;
        pixel_data[133][173] = 0;
        pixel_data[133][174] = 0;
        pixel_data[133][175] = 0;
        pixel_data[133][176] = 0;
        pixel_data[133][177] = 0;
        pixel_data[133][178] = 0;
        pixel_data[133][179] = 0;
        pixel_data[133][180] = 0;
        pixel_data[133][181] = 0;
        pixel_data[133][182] = 0;
        pixel_data[133][183] = 0;
        pixel_data[133][184] = 0;
        pixel_data[133][185] = 0;
        pixel_data[133][186] = 0;
        pixel_data[133][187] = 0;
        pixel_data[133][188] = 0;
        pixel_data[133][189] = 0;
        pixel_data[133][190] = 0;
        pixel_data[133][191] = 0;
        pixel_data[133][192] = 0;
        pixel_data[133][193] = 0;
        pixel_data[133][194] = 0;
        pixel_data[133][195] = 0;
        pixel_data[133][196] = 0;
        pixel_data[133][197] = 0;
        pixel_data[133][198] = 0;
        pixel_data[133][199] = 0; // y=133
        pixel_data[134][0] = 0;
        pixel_data[134][1] = 0;
        pixel_data[134][2] = 0;
        pixel_data[134][3] = 0;
        pixel_data[134][4] = 0;
        pixel_data[134][5] = 0;
        pixel_data[134][6] = 0;
        pixel_data[134][7] = 0;
        pixel_data[134][8] = 0;
        pixel_data[134][9] = 0;
        pixel_data[134][10] = 0;
        pixel_data[134][11] = 0;
        pixel_data[134][12] = 0;
        pixel_data[134][13] = 0;
        pixel_data[134][14] = 0;
        pixel_data[134][15] = 0;
        pixel_data[134][16] = 0;
        pixel_data[134][17] = 0;
        pixel_data[134][18] = 0;
        pixel_data[134][19] = 0;
        pixel_data[134][20] = 0;
        pixel_data[134][21] = 0;
        pixel_data[134][22] = 0;
        pixel_data[134][23] = 0;
        pixel_data[134][24] = 0;
        pixel_data[134][25] = 0;
        pixel_data[134][26] = 0;
        pixel_data[134][27] = 0;
        pixel_data[134][28] = 0;
        pixel_data[134][29] = 0;
        pixel_data[134][30] = 0;
        pixel_data[134][31] = 0;
        pixel_data[134][32] = 0;
        pixel_data[134][33] = 0;
        pixel_data[134][34] = 0;
        pixel_data[134][35] = 0;
        pixel_data[134][36] = 0;
        pixel_data[134][37] = 0;
        pixel_data[134][38] = 0;
        pixel_data[134][39] = 0;
        pixel_data[134][40] = 0;
        pixel_data[134][41] = 0;
        pixel_data[134][42] = 0;
        pixel_data[134][43] = 0;
        pixel_data[134][44] = 0;
        pixel_data[134][45] = 0;
        pixel_data[134][46] = 0;
        pixel_data[134][47] = 0;
        pixel_data[134][48] = 0;
        pixel_data[134][49] = 0;
        pixel_data[134][50] = 0;
        pixel_data[134][51] = 0;
        pixel_data[134][52] = 0;
        pixel_data[134][53] = 0;
        pixel_data[134][54] = 0;
        pixel_data[134][55] = 0;
        pixel_data[134][56] = 0;
        pixel_data[134][57] = 0;
        pixel_data[134][58] = 0;
        pixel_data[134][59] = 0;
        pixel_data[134][60] = 0;
        pixel_data[134][61] = 0;
        pixel_data[134][62] = 0;
        pixel_data[134][63] = 0;
        pixel_data[134][64] = 0;
        pixel_data[134][65] = 0;
        pixel_data[134][66] = 0;
        pixel_data[134][67] = 0;
        pixel_data[134][68] = 0;
        pixel_data[134][69] = 0;
        pixel_data[134][70] = 0;
        pixel_data[134][71] = 0;
        pixel_data[134][72] = 0;
        pixel_data[134][73] = 0;
        pixel_data[134][74] = 0;
        pixel_data[134][75] = 0;
        pixel_data[134][76] = 0;
        pixel_data[134][77] = 0;
        pixel_data[134][78] = 0;
        pixel_data[134][79] = 0;
        pixel_data[134][80] = 0;
        pixel_data[134][81] = 0;
        pixel_data[134][82] = 0;
        pixel_data[134][83] = 0;
        pixel_data[134][84] = 0;
        pixel_data[134][85] = 0;
        pixel_data[134][86] = 0;
        pixel_data[134][87] = 0;
        pixel_data[134][88] = 0;
        pixel_data[134][89] = 0;
        pixel_data[134][90] = 0;
        pixel_data[134][91] = 0;
        pixel_data[134][92] = 0;
        pixel_data[134][93] = 0;
        pixel_data[134][94] = 0;
        pixel_data[134][95] = 0;
        pixel_data[134][96] = 0;
        pixel_data[134][97] = 0;
        pixel_data[134][98] = 0;
        pixel_data[134][99] = 0;
        pixel_data[134][100] = 0;
        pixel_data[134][101] = 0;
        pixel_data[134][102] = 0;
        pixel_data[134][103] = 0;
        pixel_data[134][104] = 0;
        pixel_data[134][105] = 0;
        pixel_data[134][106] = 0;
        pixel_data[134][107] = 0;
        pixel_data[134][108] = 0;
        pixel_data[134][109] = 0;
        pixel_data[134][110] = 0;
        pixel_data[134][111] = 0;
        pixel_data[134][112] = 0;
        pixel_data[134][113] = 0;
        pixel_data[134][114] = 0;
        pixel_data[134][115] = 0;
        pixel_data[134][116] = 0;
        pixel_data[134][117] = 0;
        pixel_data[134][118] = 0;
        pixel_data[134][119] = 0;
        pixel_data[134][120] = 0;
        pixel_data[134][121] = 0;
        pixel_data[134][122] = 0;
        pixel_data[134][123] = 0;
        pixel_data[134][124] = 0;
        pixel_data[134][125] = 0;
        pixel_data[134][126] = 0;
        pixel_data[134][127] = 0;
        pixel_data[134][128] = 0;
        pixel_data[134][129] = 0;
        pixel_data[134][130] = 0;
        pixel_data[134][131] = 0;
        pixel_data[134][132] = 0;
        pixel_data[134][133] = 0;
        pixel_data[134][134] = 0;
        pixel_data[134][135] = 0;
        pixel_data[134][136] = 0;
        pixel_data[134][137] = 0;
        pixel_data[134][138] = 0;
        pixel_data[134][139] = 0;
        pixel_data[134][140] = 0;
        pixel_data[134][141] = 0;
        pixel_data[134][142] = 0;
        pixel_data[134][143] = 0;
        pixel_data[134][144] = 0;
        pixel_data[134][145] = 0;
        pixel_data[134][146] = 0;
        pixel_data[134][147] = 0;
        pixel_data[134][148] = 0;
        pixel_data[134][149] = 0;
        pixel_data[134][150] = 0;
        pixel_data[134][151] = 0;
        pixel_data[134][152] = 0;
        pixel_data[134][153] = 0;
        pixel_data[134][154] = 0;
        pixel_data[134][155] = 0;
        pixel_data[134][156] = 0;
        pixel_data[134][157] = 0;
        pixel_data[134][158] = 0;
        pixel_data[134][159] = 0;
        pixel_data[134][160] = 0;
        pixel_data[134][161] = 0;
        pixel_data[134][162] = 0;
        pixel_data[134][163] = 0;
        pixel_data[134][164] = 0;
        pixel_data[134][165] = 0;
        pixel_data[134][166] = 0;
        pixel_data[134][167] = 0;
        pixel_data[134][168] = 0;
        pixel_data[134][169] = 0;
        pixel_data[134][170] = 0;
        pixel_data[134][171] = 0;
        pixel_data[134][172] = 0;
        pixel_data[134][173] = 0;
        pixel_data[134][174] = 0;
        pixel_data[134][175] = 0;
        pixel_data[134][176] = 0;
        pixel_data[134][177] = 0;
        pixel_data[134][178] = 0;
        pixel_data[134][179] = 0;
        pixel_data[134][180] = 0;
        pixel_data[134][181] = 0;
        pixel_data[134][182] = 0;
        pixel_data[134][183] = 0;
        pixel_data[134][184] = 0;
        pixel_data[134][185] = 0;
        pixel_data[134][186] = 0;
        pixel_data[134][187] = 0;
        pixel_data[134][188] = 0;
        pixel_data[134][189] = 0;
        pixel_data[134][190] = 0;
        pixel_data[134][191] = 0;
        pixel_data[134][192] = 0;
        pixel_data[134][193] = 0;
        pixel_data[134][194] = 0;
        pixel_data[134][195] = 0;
        pixel_data[134][196] = 0;
        pixel_data[134][197] = 0;
        pixel_data[134][198] = 0;
        pixel_data[134][199] = 0; // y=134
        pixel_data[135][0] = 0;
        pixel_data[135][1] = 0;
        pixel_data[135][2] = 0;
        pixel_data[135][3] = 0;
        pixel_data[135][4] = 0;
        pixel_data[135][5] = 0;
        pixel_data[135][6] = 0;
        pixel_data[135][7] = 0;
        pixel_data[135][8] = 0;
        pixel_data[135][9] = 0;
        pixel_data[135][10] = 0;
        pixel_data[135][11] = 0;
        pixel_data[135][12] = 0;
        pixel_data[135][13] = 0;
        pixel_data[135][14] = 0;
        pixel_data[135][15] = 0;
        pixel_data[135][16] = 0;
        pixel_data[135][17] = 0;
        pixel_data[135][18] = 0;
        pixel_data[135][19] = 0;
        pixel_data[135][20] = 0;
        pixel_data[135][21] = 0;
        pixel_data[135][22] = 0;
        pixel_data[135][23] = 0;
        pixel_data[135][24] = 0;
        pixel_data[135][25] = 0;
        pixel_data[135][26] = 0;
        pixel_data[135][27] = 0;
        pixel_data[135][28] = 0;
        pixel_data[135][29] = 0;
        pixel_data[135][30] = 0;
        pixel_data[135][31] = 0;
        pixel_data[135][32] = 0;
        pixel_data[135][33] = 0;
        pixel_data[135][34] = 0;
        pixel_data[135][35] = 0;
        pixel_data[135][36] = 0;
        pixel_data[135][37] = 0;
        pixel_data[135][38] = 0;
        pixel_data[135][39] = 0;
        pixel_data[135][40] = 0;
        pixel_data[135][41] = 0;
        pixel_data[135][42] = 0;
        pixel_data[135][43] = 0;
        pixel_data[135][44] = 0;
        pixel_data[135][45] = 0;
        pixel_data[135][46] = 0;
        pixel_data[135][47] = 0;
        pixel_data[135][48] = 0;
        pixel_data[135][49] = 0;
        pixel_data[135][50] = 0;
        pixel_data[135][51] = 0;
        pixel_data[135][52] = 0;
        pixel_data[135][53] = 0;
        pixel_data[135][54] = 0;
        pixel_data[135][55] = 0;
        pixel_data[135][56] = 0;
        pixel_data[135][57] = 0;
        pixel_data[135][58] = 0;
        pixel_data[135][59] = 0;
        pixel_data[135][60] = 0;
        pixel_data[135][61] = 0;
        pixel_data[135][62] = 0;
        pixel_data[135][63] = 0;
        pixel_data[135][64] = 0;
        pixel_data[135][65] = 0;
        pixel_data[135][66] = 0;
        pixel_data[135][67] = 0;
        pixel_data[135][68] = 0;
        pixel_data[135][69] = 0;
        pixel_data[135][70] = 0;
        pixel_data[135][71] = 0;
        pixel_data[135][72] = 0;
        pixel_data[135][73] = 0;
        pixel_data[135][74] = 0;
        pixel_data[135][75] = 0;
        pixel_data[135][76] = 0;
        pixel_data[135][77] = 0;
        pixel_data[135][78] = 0;
        pixel_data[135][79] = 0;
        pixel_data[135][80] = 0;
        pixel_data[135][81] = 0;
        pixel_data[135][82] = 0;
        pixel_data[135][83] = 0;
        pixel_data[135][84] = 0;
        pixel_data[135][85] = 0;
        pixel_data[135][86] = 0;
        pixel_data[135][87] = 0;
        pixel_data[135][88] = 0;
        pixel_data[135][89] = 0;
        pixel_data[135][90] = 0;
        pixel_data[135][91] = 0;
        pixel_data[135][92] = 0;
        pixel_data[135][93] = 0;
        pixel_data[135][94] = 0;
        pixel_data[135][95] = 0;
        pixel_data[135][96] = 0;
        pixel_data[135][97] = 0;
        pixel_data[135][98] = 0;
        pixel_data[135][99] = 0;
        pixel_data[135][100] = 0;
        pixel_data[135][101] = 0;
        pixel_data[135][102] = 0;
        pixel_data[135][103] = 0;
        pixel_data[135][104] = 0;
        pixel_data[135][105] = 0;
        pixel_data[135][106] = 0;
        pixel_data[135][107] = 0;
        pixel_data[135][108] = 0;
        pixel_data[135][109] = 0;
        pixel_data[135][110] = 0;
        pixel_data[135][111] = 0;
        pixel_data[135][112] = 0;
        pixel_data[135][113] = 0;
        pixel_data[135][114] = 0;
        pixel_data[135][115] = 0;
        pixel_data[135][116] = 0;
        pixel_data[135][117] = 0;
        pixel_data[135][118] = 0;
        pixel_data[135][119] = 0;
        pixel_data[135][120] = 0;
        pixel_data[135][121] = 0;
        pixel_data[135][122] = 0;
        pixel_data[135][123] = 0;
        pixel_data[135][124] = 0;
        pixel_data[135][125] = 0;
        pixel_data[135][126] = 0;
        pixel_data[135][127] = 0;
        pixel_data[135][128] = 0;
        pixel_data[135][129] = 0;
        pixel_data[135][130] = 0;
        pixel_data[135][131] = 0;
        pixel_data[135][132] = 0;
        pixel_data[135][133] = 0;
        pixel_data[135][134] = 0;
        pixel_data[135][135] = 0;
        pixel_data[135][136] = 0;
        pixel_data[135][137] = 0;
        pixel_data[135][138] = 0;
        pixel_data[135][139] = 0;
        pixel_data[135][140] = 0;
        pixel_data[135][141] = 0;
        pixel_data[135][142] = 0;
        pixel_data[135][143] = 0;
        pixel_data[135][144] = 0;
        pixel_data[135][145] = 0;
        pixel_data[135][146] = 0;
        pixel_data[135][147] = 0;
        pixel_data[135][148] = 0;
        pixel_data[135][149] = 0;
        pixel_data[135][150] = 0;
        pixel_data[135][151] = 0;
        pixel_data[135][152] = 0;
        pixel_data[135][153] = 0;
        pixel_data[135][154] = 0;
        pixel_data[135][155] = 0;
        pixel_data[135][156] = 0;
        pixel_data[135][157] = 0;
        pixel_data[135][158] = 0;
        pixel_data[135][159] = 0;
        pixel_data[135][160] = 0;
        pixel_data[135][161] = 0;
        pixel_data[135][162] = 0;
        pixel_data[135][163] = 0;
        pixel_data[135][164] = 0;
        pixel_data[135][165] = 0;
        pixel_data[135][166] = 0;
        pixel_data[135][167] = 0;
        pixel_data[135][168] = 0;
        pixel_data[135][169] = 0;
        pixel_data[135][170] = 0;
        pixel_data[135][171] = 0;
        pixel_data[135][172] = 0;
        pixel_data[135][173] = 0;
        pixel_data[135][174] = 0;
        pixel_data[135][175] = 0;
        pixel_data[135][176] = 0;
        pixel_data[135][177] = 0;
        pixel_data[135][178] = 0;
        pixel_data[135][179] = 0;
        pixel_data[135][180] = 0;
        pixel_data[135][181] = 0;
        pixel_data[135][182] = 0;
        pixel_data[135][183] = 0;
        pixel_data[135][184] = 0;
        pixel_data[135][185] = 0;
        pixel_data[135][186] = 0;
        pixel_data[135][187] = 0;
        pixel_data[135][188] = 0;
        pixel_data[135][189] = 0;
        pixel_data[135][190] = 0;
        pixel_data[135][191] = 0;
        pixel_data[135][192] = 0;
        pixel_data[135][193] = 0;
        pixel_data[135][194] = 0;
        pixel_data[135][195] = 0;
        pixel_data[135][196] = 0;
        pixel_data[135][197] = 0;
        pixel_data[135][198] = 0;
        pixel_data[135][199] = 0; // y=135
        pixel_data[136][0] = 0;
        pixel_data[136][1] = 0;
        pixel_data[136][2] = 0;
        pixel_data[136][3] = 0;
        pixel_data[136][4] = 0;
        pixel_data[136][5] = 0;
        pixel_data[136][6] = 0;
        pixel_data[136][7] = 0;
        pixel_data[136][8] = 0;
        pixel_data[136][9] = 0;
        pixel_data[136][10] = 0;
        pixel_data[136][11] = 0;
        pixel_data[136][12] = 0;
        pixel_data[136][13] = 0;
        pixel_data[136][14] = 0;
        pixel_data[136][15] = 0;
        pixel_data[136][16] = 0;
        pixel_data[136][17] = 0;
        pixel_data[136][18] = 0;
        pixel_data[136][19] = 0;
        pixel_data[136][20] = 0;
        pixel_data[136][21] = 0;
        pixel_data[136][22] = 0;
        pixel_data[136][23] = 0;
        pixel_data[136][24] = 0;
        pixel_data[136][25] = 0;
        pixel_data[136][26] = 0;
        pixel_data[136][27] = 0;
        pixel_data[136][28] = 0;
        pixel_data[136][29] = 0;
        pixel_data[136][30] = 0;
        pixel_data[136][31] = 0;
        pixel_data[136][32] = 0;
        pixel_data[136][33] = 0;
        pixel_data[136][34] = 0;
        pixel_data[136][35] = 0;
        pixel_data[136][36] = 0;
        pixel_data[136][37] = 0;
        pixel_data[136][38] = 0;
        pixel_data[136][39] = 0;
        pixel_data[136][40] = 0;
        pixel_data[136][41] = 0;
        pixel_data[136][42] = 0;
        pixel_data[136][43] = 0;
        pixel_data[136][44] = 0;
        pixel_data[136][45] = 0;
        pixel_data[136][46] = 0;
        pixel_data[136][47] = 0;
        pixel_data[136][48] = 0;
        pixel_data[136][49] = 0;
        pixel_data[136][50] = 0;
        pixel_data[136][51] = 0;
        pixel_data[136][52] = 0;
        pixel_data[136][53] = 0;
        pixel_data[136][54] = 0;
        pixel_data[136][55] = 0;
        pixel_data[136][56] = 0;
        pixel_data[136][57] = 0;
        pixel_data[136][58] = 0;
        pixel_data[136][59] = 0;
        pixel_data[136][60] = 0;
        pixel_data[136][61] = 0;
        pixel_data[136][62] = 0;
        pixel_data[136][63] = 0;
        pixel_data[136][64] = 0;
        pixel_data[136][65] = 0;
        pixel_data[136][66] = 0;
        pixel_data[136][67] = 0;
        pixel_data[136][68] = 0;
        pixel_data[136][69] = 0;
        pixel_data[136][70] = 0;
        pixel_data[136][71] = 0;
        pixel_data[136][72] = 0;
        pixel_data[136][73] = 0;
        pixel_data[136][74] = 0;
        pixel_data[136][75] = 0;
        pixel_data[136][76] = 0;
        pixel_data[136][77] = 0;
        pixel_data[136][78] = 0;
        pixel_data[136][79] = 0;
        pixel_data[136][80] = 0;
        pixel_data[136][81] = 0;
        pixel_data[136][82] = 0;
        pixel_data[136][83] = 0;
        pixel_data[136][84] = 0;
        pixel_data[136][85] = 0;
        pixel_data[136][86] = 0;
        pixel_data[136][87] = 0;
        pixel_data[136][88] = 0;
        pixel_data[136][89] = 0;
        pixel_data[136][90] = 0;
        pixel_data[136][91] = 0;
        pixel_data[136][92] = 0;
        pixel_data[136][93] = 0;
        pixel_data[136][94] = 0;
        pixel_data[136][95] = 0;
        pixel_data[136][96] = 0;
        pixel_data[136][97] = 0;
        pixel_data[136][98] = 0;
        pixel_data[136][99] = 0;
        pixel_data[136][100] = 0;
        pixel_data[136][101] = 0;
        pixel_data[136][102] = 0;
        pixel_data[136][103] = 0;
        pixel_data[136][104] = 0;
        pixel_data[136][105] = 0;
        pixel_data[136][106] = 0;
        pixel_data[136][107] = 0;
        pixel_data[136][108] = 0;
        pixel_data[136][109] = 0;
        pixel_data[136][110] = 0;
        pixel_data[136][111] = 0;
        pixel_data[136][112] = 0;
        pixel_data[136][113] = 0;
        pixel_data[136][114] = 0;
        pixel_data[136][115] = 0;
        pixel_data[136][116] = 0;
        pixel_data[136][117] = 0;
        pixel_data[136][118] = 0;
        pixel_data[136][119] = 0;
        pixel_data[136][120] = 0;
        pixel_data[136][121] = 0;
        pixel_data[136][122] = 0;
        pixel_data[136][123] = 0;
        pixel_data[136][124] = 0;
        pixel_data[136][125] = 0;
        pixel_data[136][126] = 0;
        pixel_data[136][127] = 0;
        pixel_data[136][128] = 0;
        pixel_data[136][129] = 0;
        pixel_data[136][130] = 0;
        pixel_data[136][131] = 0;
        pixel_data[136][132] = 0;
        pixel_data[136][133] = 0;
        pixel_data[136][134] = 0;
        pixel_data[136][135] = 0;
        pixel_data[136][136] = 0;
        pixel_data[136][137] = 0;
        pixel_data[136][138] = 0;
        pixel_data[136][139] = 0;
        pixel_data[136][140] = 0;
        pixel_data[136][141] = 0;
        pixel_data[136][142] = 0;
        pixel_data[136][143] = 0;
        pixel_data[136][144] = 0;
        pixel_data[136][145] = 0;
        pixel_data[136][146] = 0;
        pixel_data[136][147] = 0;
        pixel_data[136][148] = 0;
        pixel_data[136][149] = 0;
        pixel_data[136][150] = 0;
        pixel_data[136][151] = 0;
        pixel_data[136][152] = 0;
        pixel_data[136][153] = 0;
        pixel_data[136][154] = 0;
        pixel_data[136][155] = 0;
        pixel_data[136][156] = 0;
        pixel_data[136][157] = 0;
        pixel_data[136][158] = 0;
        pixel_data[136][159] = 0;
        pixel_data[136][160] = 0;
        pixel_data[136][161] = 0;
        pixel_data[136][162] = 0;
        pixel_data[136][163] = 0;
        pixel_data[136][164] = 0;
        pixel_data[136][165] = 0;
        pixel_data[136][166] = 0;
        pixel_data[136][167] = 0;
        pixel_data[136][168] = 0;
        pixel_data[136][169] = 0;
        pixel_data[136][170] = 0;
        pixel_data[136][171] = 0;
        pixel_data[136][172] = 0;
        pixel_data[136][173] = 0;
        pixel_data[136][174] = 0;
        pixel_data[136][175] = 0;
        pixel_data[136][176] = 0;
        pixel_data[136][177] = 0;
        pixel_data[136][178] = 0;
        pixel_data[136][179] = 0;
        pixel_data[136][180] = 0;
        pixel_data[136][181] = 0;
        pixel_data[136][182] = 0;
        pixel_data[136][183] = 0;
        pixel_data[136][184] = 0;
        pixel_data[136][185] = 0;
        pixel_data[136][186] = 0;
        pixel_data[136][187] = 0;
        pixel_data[136][188] = 0;
        pixel_data[136][189] = 0;
        pixel_data[136][190] = 0;
        pixel_data[136][191] = 0;
        pixel_data[136][192] = 0;
        pixel_data[136][193] = 0;
        pixel_data[136][194] = 0;
        pixel_data[136][195] = 0;
        pixel_data[136][196] = 0;
        pixel_data[136][197] = 0;
        pixel_data[136][198] = 0;
        pixel_data[136][199] = 0; // y=136
        pixel_data[137][0] = 0;
        pixel_data[137][1] = 0;
        pixel_data[137][2] = 0;
        pixel_data[137][3] = 0;
        pixel_data[137][4] = 0;
        pixel_data[137][5] = 0;
        pixel_data[137][6] = 0;
        pixel_data[137][7] = 0;
        pixel_data[137][8] = 0;
        pixel_data[137][9] = 0;
        pixel_data[137][10] = 0;
        pixel_data[137][11] = 0;
        pixel_data[137][12] = 0;
        pixel_data[137][13] = 0;
        pixel_data[137][14] = 0;
        pixel_data[137][15] = 0;
        pixel_data[137][16] = 0;
        pixel_data[137][17] = 0;
        pixel_data[137][18] = 0;
        pixel_data[137][19] = 0;
        pixel_data[137][20] = 0;
        pixel_data[137][21] = 0;
        pixel_data[137][22] = 0;
        pixel_data[137][23] = 0;
        pixel_data[137][24] = 0;
        pixel_data[137][25] = 0;
        pixel_data[137][26] = 0;
        pixel_data[137][27] = 0;
        pixel_data[137][28] = 0;
        pixel_data[137][29] = 0;
        pixel_data[137][30] = 0;
        pixel_data[137][31] = 0;
        pixel_data[137][32] = 0;
        pixel_data[137][33] = 0;
        pixel_data[137][34] = 0;
        pixel_data[137][35] = 0;
        pixel_data[137][36] = 0;
        pixel_data[137][37] = 0;
        pixel_data[137][38] = 0;
        pixel_data[137][39] = 0;
        pixel_data[137][40] = 0;
        pixel_data[137][41] = 0;
        pixel_data[137][42] = 0;
        pixel_data[137][43] = 0;
        pixel_data[137][44] = 0;
        pixel_data[137][45] = 0;
        pixel_data[137][46] = 0;
        pixel_data[137][47] = 0;
        pixel_data[137][48] = 0;
        pixel_data[137][49] = 0;
        pixel_data[137][50] = 0;
        pixel_data[137][51] = 0;
        pixel_data[137][52] = 0;
        pixel_data[137][53] = 0;
        pixel_data[137][54] = 0;
        pixel_data[137][55] = 0;
        pixel_data[137][56] = 0;
        pixel_data[137][57] = 0;
        pixel_data[137][58] = 0;
        pixel_data[137][59] = 0;
        pixel_data[137][60] = 0;
        pixel_data[137][61] = 0;
        pixel_data[137][62] = 0;
        pixel_data[137][63] = 0;
        pixel_data[137][64] = 0;
        pixel_data[137][65] = 0;
        pixel_data[137][66] = 0;
        pixel_data[137][67] = 0;
        pixel_data[137][68] = 0;
        pixel_data[137][69] = 0;
        pixel_data[137][70] = 0;
        pixel_data[137][71] = 0;
        pixel_data[137][72] = 0;
        pixel_data[137][73] = 0;
        pixel_data[137][74] = 0;
        pixel_data[137][75] = 0;
        pixel_data[137][76] = 0;
        pixel_data[137][77] = 0;
        pixel_data[137][78] = 0;
        pixel_data[137][79] = 0;
        pixel_data[137][80] = 0;
        pixel_data[137][81] = 0;
        pixel_data[137][82] = 0;
        pixel_data[137][83] = 0;
        pixel_data[137][84] = 0;
        pixel_data[137][85] = 0;
        pixel_data[137][86] = 0;
        pixel_data[137][87] = 0;
        pixel_data[137][88] = 0;
        pixel_data[137][89] = 0;
        pixel_data[137][90] = 0;
        pixel_data[137][91] = 0;
        pixel_data[137][92] = 0;
        pixel_data[137][93] = 0;
        pixel_data[137][94] = 0;
        pixel_data[137][95] = 0;
        pixel_data[137][96] = 0;
        pixel_data[137][97] = 0;
        pixel_data[137][98] = 0;
        pixel_data[137][99] = 0;
        pixel_data[137][100] = 0;
        pixel_data[137][101] = 0;
        pixel_data[137][102] = 0;
        pixel_data[137][103] = 0;
        pixel_data[137][104] = 0;
        pixel_data[137][105] = 0;
        pixel_data[137][106] = 0;
        pixel_data[137][107] = 0;
        pixel_data[137][108] = 0;
        pixel_data[137][109] = 0;
        pixel_data[137][110] = 0;
        pixel_data[137][111] = 0;
        pixel_data[137][112] = 0;
        pixel_data[137][113] = 0;
        pixel_data[137][114] = 0;
        pixel_data[137][115] = 0;
        pixel_data[137][116] = 0;
        pixel_data[137][117] = 0;
        pixel_data[137][118] = 0;
        pixel_data[137][119] = 0;
        pixel_data[137][120] = 0;
        pixel_data[137][121] = 0;
        pixel_data[137][122] = 0;
        pixel_data[137][123] = 0;
        pixel_data[137][124] = 0;
        pixel_data[137][125] = 0;
        pixel_data[137][126] = 0;
        pixel_data[137][127] = 0;
        pixel_data[137][128] = 0;
        pixel_data[137][129] = 0;
        pixel_data[137][130] = 0;
        pixel_data[137][131] = 0;
        pixel_data[137][132] = 0;
        pixel_data[137][133] = 0;
        pixel_data[137][134] = 0;
        pixel_data[137][135] = 0;
        pixel_data[137][136] = 0;
        pixel_data[137][137] = 0;
        pixel_data[137][138] = 0;
        pixel_data[137][139] = 0;
        pixel_data[137][140] = 0;
        pixel_data[137][141] = 0;
        pixel_data[137][142] = 0;
        pixel_data[137][143] = 0;
        pixel_data[137][144] = 0;
        pixel_data[137][145] = 0;
        pixel_data[137][146] = 0;
        pixel_data[137][147] = 0;
        pixel_data[137][148] = 0;
        pixel_data[137][149] = 0;
        pixel_data[137][150] = 0;
        pixel_data[137][151] = 0;
        pixel_data[137][152] = 0;
        pixel_data[137][153] = 0;
        pixel_data[137][154] = 0;
        pixel_data[137][155] = 0;
        pixel_data[137][156] = 0;
        pixel_data[137][157] = 0;
        pixel_data[137][158] = 0;
        pixel_data[137][159] = 0;
        pixel_data[137][160] = 0;
        pixel_data[137][161] = 0;
        pixel_data[137][162] = 0;
        pixel_data[137][163] = 0;
        pixel_data[137][164] = 0;
        pixel_data[137][165] = 0;
        pixel_data[137][166] = 0;
        pixel_data[137][167] = 0;
        pixel_data[137][168] = 0;
        pixel_data[137][169] = 0;
        pixel_data[137][170] = 0;
        pixel_data[137][171] = 0;
        pixel_data[137][172] = 0;
        pixel_data[137][173] = 0;
        pixel_data[137][174] = 0;
        pixel_data[137][175] = 0;
        pixel_data[137][176] = 0;
        pixel_data[137][177] = 0;
        pixel_data[137][178] = 0;
        pixel_data[137][179] = 0;
        pixel_data[137][180] = 0;
        pixel_data[137][181] = 0;
        pixel_data[137][182] = 0;
        pixel_data[137][183] = 0;
        pixel_data[137][184] = 0;
        pixel_data[137][185] = 0;
        pixel_data[137][186] = 0;
        pixel_data[137][187] = 0;
        pixel_data[137][188] = 0;
        pixel_data[137][189] = 0;
        pixel_data[137][190] = 0;
        pixel_data[137][191] = 0;
        pixel_data[137][192] = 0;
        pixel_data[137][193] = 0;
        pixel_data[137][194] = 0;
        pixel_data[137][195] = 0;
        pixel_data[137][196] = 0;
        pixel_data[137][197] = 0;
        pixel_data[137][198] = 0;
        pixel_data[137][199] = 0; // y=137
        pixel_data[138][0] = 0;
        pixel_data[138][1] = 0;
        pixel_data[138][2] = 0;
        pixel_data[138][3] = 0;
        pixel_data[138][4] = 0;
        pixel_data[138][5] = 0;
        pixel_data[138][6] = 0;
        pixel_data[138][7] = 0;
        pixel_data[138][8] = 0;
        pixel_data[138][9] = 0;
        pixel_data[138][10] = 0;
        pixel_data[138][11] = 0;
        pixel_data[138][12] = 0;
        pixel_data[138][13] = 0;
        pixel_data[138][14] = 0;
        pixel_data[138][15] = 0;
        pixel_data[138][16] = 0;
        pixel_data[138][17] = 0;
        pixel_data[138][18] = 0;
        pixel_data[138][19] = 0;
        pixel_data[138][20] = 0;
        pixel_data[138][21] = 0;
        pixel_data[138][22] = 0;
        pixel_data[138][23] = 0;
        pixel_data[138][24] = 0;
        pixel_data[138][25] = 0;
        pixel_data[138][26] = 0;
        pixel_data[138][27] = 0;
        pixel_data[138][28] = 0;
        pixel_data[138][29] = 0;
        pixel_data[138][30] = 0;
        pixel_data[138][31] = 0;
        pixel_data[138][32] = 0;
        pixel_data[138][33] = 0;
        pixel_data[138][34] = 0;
        pixel_data[138][35] = 0;
        pixel_data[138][36] = 0;
        pixel_data[138][37] = 0;
        pixel_data[138][38] = 0;
        pixel_data[138][39] = 0;
        pixel_data[138][40] = 0;
        pixel_data[138][41] = 0;
        pixel_data[138][42] = 0;
        pixel_data[138][43] = 0;
        pixel_data[138][44] = 0;
        pixel_data[138][45] = 0;
        pixel_data[138][46] = 0;
        pixel_data[138][47] = 0;
        pixel_data[138][48] = 0;
        pixel_data[138][49] = 0;
        pixel_data[138][50] = 0;
        pixel_data[138][51] = 0;
        pixel_data[138][52] = 0;
        pixel_data[138][53] = 0;
        pixel_data[138][54] = 0;
        pixel_data[138][55] = 0;
        pixel_data[138][56] = 0;
        pixel_data[138][57] = 0;
        pixel_data[138][58] = 0;
        pixel_data[138][59] = 0;
        pixel_data[138][60] = 0;
        pixel_data[138][61] = 0;
        pixel_data[138][62] = 0;
        pixel_data[138][63] = 0;
        pixel_data[138][64] = 0;
        pixel_data[138][65] = 0;
        pixel_data[138][66] = 0;
        pixel_data[138][67] = 0;
        pixel_data[138][68] = 0;
        pixel_data[138][69] = 0;
        pixel_data[138][70] = 0;
        pixel_data[138][71] = 0;
        pixel_data[138][72] = 0;
        pixel_data[138][73] = 0;
        pixel_data[138][74] = 0;
        pixel_data[138][75] = 0;
        pixel_data[138][76] = 0;
        pixel_data[138][77] = 0;
        pixel_data[138][78] = 0;
        pixel_data[138][79] = 0;
        pixel_data[138][80] = 0;
        pixel_data[138][81] = 0;
        pixel_data[138][82] = 0;
        pixel_data[138][83] = 0;
        pixel_data[138][84] = 0;
        pixel_data[138][85] = 0;
        pixel_data[138][86] = 0;
        pixel_data[138][87] = 0;
        pixel_data[138][88] = 0;
        pixel_data[138][89] = 0;
        pixel_data[138][90] = 0;
        pixel_data[138][91] = 0;
        pixel_data[138][92] = 0;
        pixel_data[138][93] = 0;
        pixel_data[138][94] = 0;
        pixel_data[138][95] = 0;
        pixel_data[138][96] = 0;
        pixel_data[138][97] = 0;
        pixel_data[138][98] = 0;
        pixel_data[138][99] = 0;
        pixel_data[138][100] = 0;
        pixel_data[138][101] = 0;
        pixel_data[138][102] = 0;
        pixel_data[138][103] = 0;
        pixel_data[138][104] = 0;
        pixel_data[138][105] = 0;
        pixel_data[138][106] = 0;
        pixel_data[138][107] = 0;
        pixel_data[138][108] = 0;
        pixel_data[138][109] = 0;
        pixel_data[138][110] = 0;
        pixel_data[138][111] = 0;
        pixel_data[138][112] = 0;
        pixel_data[138][113] = 0;
        pixel_data[138][114] = 0;
        pixel_data[138][115] = 0;
        pixel_data[138][116] = 0;
        pixel_data[138][117] = 0;
        pixel_data[138][118] = 0;
        pixel_data[138][119] = 0;
        pixel_data[138][120] = 0;
        pixel_data[138][121] = 0;
        pixel_data[138][122] = 0;
        pixel_data[138][123] = 0;
        pixel_data[138][124] = 0;
        pixel_data[138][125] = 0;
        pixel_data[138][126] = 0;
        pixel_data[138][127] = 0;
        pixel_data[138][128] = 0;
        pixel_data[138][129] = 0;
        pixel_data[138][130] = 0;
        pixel_data[138][131] = 0;
        pixel_data[138][132] = 0;
        pixel_data[138][133] = 0;
        pixel_data[138][134] = 0;
        pixel_data[138][135] = 0;
        pixel_data[138][136] = 0;
        pixel_data[138][137] = 0;
        pixel_data[138][138] = 0;
        pixel_data[138][139] = 0;
        pixel_data[138][140] = 0;
        pixel_data[138][141] = 0;
        pixel_data[138][142] = 0;
        pixel_data[138][143] = 0;
        pixel_data[138][144] = 0;
        pixel_data[138][145] = 0;
        pixel_data[138][146] = 0;
        pixel_data[138][147] = 0;
        pixel_data[138][148] = 0;
        pixel_data[138][149] = 0;
        pixel_data[138][150] = 0;
        pixel_data[138][151] = 0;
        pixel_data[138][152] = 0;
        pixel_data[138][153] = 0;
        pixel_data[138][154] = 0;
        pixel_data[138][155] = 0;
        pixel_data[138][156] = 0;
        pixel_data[138][157] = 0;
        pixel_data[138][158] = 0;
        pixel_data[138][159] = 0;
        pixel_data[138][160] = 0;
        pixel_data[138][161] = 0;
        pixel_data[138][162] = 0;
        pixel_data[138][163] = 0;
        pixel_data[138][164] = 0;
        pixel_data[138][165] = 0;
        pixel_data[138][166] = 0;
        pixel_data[138][167] = 0;
        pixel_data[138][168] = 0;
        pixel_data[138][169] = 0;
        pixel_data[138][170] = 0;
        pixel_data[138][171] = 0;
        pixel_data[138][172] = 0;
        pixel_data[138][173] = 0;
        pixel_data[138][174] = 0;
        pixel_data[138][175] = 0;
        pixel_data[138][176] = 0;
        pixel_data[138][177] = 0;
        pixel_data[138][178] = 0;
        pixel_data[138][179] = 0;
        pixel_data[138][180] = 0;
        pixel_data[138][181] = 0;
        pixel_data[138][182] = 0;
        pixel_data[138][183] = 0;
        pixel_data[138][184] = 0;
        pixel_data[138][185] = 0;
        pixel_data[138][186] = 0;
        pixel_data[138][187] = 0;
        pixel_data[138][188] = 0;
        pixel_data[138][189] = 0;
        pixel_data[138][190] = 0;
        pixel_data[138][191] = 0;
        pixel_data[138][192] = 0;
        pixel_data[138][193] = 0;
        pixel_data[138][194] = 0;
        pixel_data[138][195] = 0;
        pixel_data[138][196] = 0;
        pixel_data[138][197] = 0;
        pixel_data[138][198] = 0;
        pixel_data[138][199] = 0; // y=138
        pixel_data[139][0] = 0;
        pixel_data[139][1] = 0;
        pixel_data[139][2] = 0;
        pixel_data[139][3] = 0;
        pixel_data[139][4] = 0;
        pixel_data[139][5] = 0;
        pixel_data[139][6] = 0;
        pixel_data[139][7] = 0;
        pixel_data[139][8] = 0;
        pixel_data[139][9] = 0;
        pixel_data[139][10] = 0;
        pixel_data[139][11] = 0;
        pixel_data[139][12] = 0;
        pixel_data[139][13] = 0;
        pixel_data[139][14] = 0;
        pixel_data[139][15] = 0;
        pixel_data[139][16] = 0;
        pixel_data[139][17] = 0;
        pixel_data[139][18] = 0;
        pixel_data[139][19] = 0;
        pixel_data[139][20] = 0;
        pixel_data[139][21] = 0;
        pixel_data[139][22] = 0;
        pixel_data[139][23] = 0;
        pixel_data[139][24] = 0;
        pixel_data[139][25] = 0;
        pixel_data[139][26] = 0;
        pixel_data[139][27] = 0;
        pixel_data[139][28] = 0;
        pixel_data[139][29] = 0;
        pixel_data[139][30] = 0;
        pixel_data[139][31] = 0;
        pixel_data[139][32] = 0;
        pixel_data[139][33] = 0;
        pixel_data[139][34] = 0;
        pixel_data[139][35] = 0;
        pixel_data[139][36] = 0;
        pixel_data[139][37] = 0;
        pixel_data[139][38] = 0;
        pixel_data[139][39] = 0;
        pixel_data[139][40] = 0;
        pixel_data[139][41] = 0;
        pixel_data[139][42] = 0;
        pixel_data[139][43] = 0;
        pixel_data[139][44] = 0;
        pixel_data[139][45] = 0;
        pixel_data[139][46] = 0;
        pixel_data[139][47] = 0;
        pixel_data[139][48] = 0;
        pixel_data[139][49] = 0;
        pixel_data[139][50] = 0;
        pixel_data[139][51] = 0;
        pixel_data[139][52] = 0;
        pixel_data[139][53] = 0;
        pixel_data[139][54] = 0;
        pixel_data[139][55] = 0;
        pixel_data[139][56] = 0;
        pixel_data[139][57] = 0;
        pixel_data[139][58] = 0;
        pixel_data[139][59] = 0;
        pixel_data[139][60] = 0;
        pixel_data[139][61] = 0;
        pixel_data[139][62] = 0;
        pixel_data[139][63] = 0;
        pixel_data[139][64] = 0;
        pixel_data[139][65] = 0;
        pixel_data[139][66] = 0;
        pixel_data[139][67] = 0;
        pixel_data[139][68] = 0;
        pixel_data[139][69] = 0;
        pixel_data[139][70] = 0;
        pixel_data[139][71] = 0;
        pixel_data[139][72] = 0;
        pixel_data[139][73] = 0;
        pixel_data[139][74] = 0;
        pixel_data[139][75] = 0;
        pixel_data[139][76] = 0;
        pixel_data[139][77] = 0;
        pixel_data[139][78] = 0;
        pixel_data[139][79] = 0;
        pixel_data[139][80] = 0;
        pixel_data[139][81] = 10;
        pixel_data[139][82] = 0;
        pixel_data[139][83] = 0;
        pixel_data[139][84] = 0;
        pixel_data[139][85] = 0;
        pixel_data[139][86] = 0;
        pixel_data[139][87] = 0;
        pixel_data[139][88] = 0;
        pixel_data[139][89] = 0;
        pixel_data[139][90] = 0;
        pixel_data[139][91] = 0;
        pixel_data[139][92] = 0;
        pixel_data[139][93] = 0;
        pixel_data[139][94] = 0;
        pixel_data[139][95] = 0;
        pixel_data[139][96] = 0;
        pixel_data[139][97] = 0;
        pixel_data[139][98] = 0;
        pixel_data[139][99] = 0;
        pixel_data[139][100] = 0;
        pixel_data[139][101] = 0;
        pixel_data[139][102] = 0;
        pixel_data[139][103] = 0;
        pixel_data[139][104] = 0;
        pixel_data[139][105] = 0;
        pixel_data[139][106] = 0;
        pixel_data[139][107] = 0;
        pixel_data[139][108] = 0;
        pixel_data[139][109] = 0;
        pixel_data[139][110] = 0;
        pixel_data[139][111] = 0;
        pixel_data[139][112] = 0;
        pixel_data[139][113] = 0;
        pixel_data[139][114] = 0;
        pixel_data[139][115] = 0;
        pixel_data[139][116] = 0;
        pixel_data[139][117] = 0;
        pixel_data[139][118] = 0;
        pixel_data[139][119] = 0;
        pixel_data[139][120] = 0;
        pixel_data[139][121] = 0;
        pixel_data[139][122] = 0;
        pixel_data[139][123] = 0;
        pixel_data[139][124] = 0;
        pixel_data[139][125] = 0;
        pixel_data[139][126] = 0;
        pixel_data[139][127] = 0;
        pixel_data[139][128] = 0;
        pixel_data[139][129] = 0;
        pixel_data[139][130] = 0;
        pixel_data[139][131] = 0;
        pixel_data[139][132] = 0;
        pixel_data[139][133] = 0;
        pixel_data[139][134] = 0;
        pixel_data[139][135] = 0;
        pixel_data[139][136] = 0;
        pixel_data[139][137] = 0;
        pixel_data[139][138] = 0;
        pixel_data[139][139] = 0;
        pixel_data[139][140] = 0;
        pixel_data[139][141] = 0;
        pixel_data[139][142] = 0;
        pixel_data[139][143] = 0;
        pixel_data[139][144] = 0;
        pixel_data[139][145] = 0;
        pixel_data[139][146] = 0;
        pixel_data[139][147] = 0;
        pixel_data[139][148] = 0;
        pixel_data[139][149] = 0;
        pixel_data[139][150] = 0;
        pixel_data[139][151] = 0;
        pixel_data[139][152] = 0;
        pixel_data[139][153] = 0;
        pixel_data[139][154] = 0;
        pixel_data[139][155] = 0;
        pixel_data[139][156] = 0;
        pixel_data[139][157] = 0;
        pixel_data[139][158] = 0;
        pixel_data[139][159] = 0;
        pixel_data[139][160] = 0;
        pixel_data[139][161] = 0;
        pixel_data[139][162] = 0;
        pixel_data[139][163] = 0;
        pixel_data[139][164] = 0;
        pixel_data[139][165] = 0;
        pixel_data[139][166] = 0;
        pixel_data[139][167] = 0;
        pixel_data[139][168] = 0;
        pixel_data[139][169] = 0;
        pixel_data[139][170] = 0;
        pixel_data[139][171] = 0;
        pixel_data[139][172] = 0;
        pixel_data[139][173] = 0;
        pixel_data[139][174] = 0;
        pixel_data[139][175] = 0;
        pixel_data[139][176] = 0;
        pixel_data[139][177] = 0;
        pixel_data[139][178] = 0;
        pixel_data[139][179] = 0;
        pixel_data[139][180] = 0;
        pixel_data[139][181] = 0;
        pixel_data[139][182] = 0;
        pixel_data[139][183] = 0;
        pixel_data[139][184] = 0;
        pixel_data[139][185] = 0;
        pixel_data[139][186] = 0;
        pixel_data[139][187] = 0;
        pixel_data[139][188] = 0;
        pixel_data[139][189] = 0;
        pixel_data[139][190] = 0;
        pixel_data[139][191] = 0;
        pixel_data[139][192] = 0;
        pixel_data[139][193] = 0;
        pixel_data[139][194] = 0;
        pixel_data[139][195] = 0;
        pixel_data[139][196] = 0;
        pixel_data[139][197] = 0;
        pixel_data[139][198] = 0;
        pixel_data[139][199] = 0; // y=139
        pixel_data[140][0] = 0;
        pixel_data[140][1] = 0;
        pixel_data[140][2] = 0;
        pixel_data[140][3] = 0;
        pixel_data[140][4] = 0;
        pixel_data[140][5] = 0;
        pixel_data[140][6] = 0;
        pixel_data[140][7] = 0;
        pixel_data[140][8] = 0;
        pixel_data[140][9] = 0;
        pixel_data[140][10] = 0;
        pixel_data[140][11] = 0;
        pixel_data[140][12] = 0;
        pixel_data[140][13] = 0;
        pixel_data[140][14] = 0;
        pixel_data[140][15] = 0;
        pixel_data[140][16] = 0;
        pixel_data[140][17] = 0;
        pixel_data[140][18] = 0;
        pixel_data[140][19] = 0;
        pixel_data[140][20] = 0;
        pixel_data[140][21] = 0;
        pixel_data[140][22] = 0;
        pixel_data[140][23] = 0;
        pixel_data[140][24] = 0;
        pixel_data[140][25] = 0;
        pixel_data[140][26] = 0;
        pixel_data[140][27] = 0;
        pixel_data[140][28] = 0;
        pixel_data[140][29] = 0;
        pixel_data[140][30] = 0;
        pixel_data[140][31] = 0;
        pixel_data[140][32] = 0;
        pixel_data[140][33] = 0;
        pixel_data[140][34] = 0;
        pixel_data[140][35] = 0;
        pixel_data[140][36] = 0;
        pixel_data[140][37] = 0;
        pixel_data[140][38] = 0;
        pixel_data[140][39] = 0;
        pixel_data[140][40] = 0;
        pixel_data[140][41] = 0;
        pixel_data[140][42] = 0;
        pixel_data[140][43] = 0;
        pixel_data[140][44] = 0;
        pixel_data[140][45] = 0;
        pixel_data[140][46] = 0;
        pixel_data[140][47] = 0;
        pixel_data[140][48] = 0;
        pixel_data[140][49] = 0;
        pixel_data[140][50] = 0;
        pixel_data[140][51] = 0;
        pixel_data[140][52] = 0;
        pixel_data[140][53] = 0;
        pixel_data[140][54] = 0;
        pixel_data[140][55] = 0;
        pixel_data[140][56] = 0;
        pixel_data[140][57] = 0;
        pixel_data[140][58] = 0;
        pixel_data[140][59] = 0;
        pixel_data[140][60] = 0;
        pixel_data[140][61] = 0;
        pixel_data[140][62] = 0;
        pixel_data[140][63] = 0;
        pixel_data[140][64] = 0;
        pixel_data[140][65] = 0;
        pixel_data[140][66] = 0;
        pixel_data[140][67] = 0;
        pixel_data[140][68] = 0;
        pixel_data[140][69] = 0;
        pixel_data[140][70] = 0;
        pixel_data[140][71] = 0;
        pixel_data[140][72] = 0;
        pixel_data[140][73] = 0;
        pixel_data[140][74] = 11;
        pixel_data[140][75] = 11;
        pixel_data[140][76] = 11;
        pixel_data[140][77] = 11;
        pixel_data[140][78] = 11;
        pixel_data[140][79] = 11;
        pixel_data[140][80] = 11;
        pixel_data[140][81] = 11;
        pixel_data[140][82] = 11;
        pixel_data[140][83] = 11;
        pixel_data[140][84] = 11;
        pixel_data[140][85] = 11;
        pixel_data[140][86] = 11;
        pixel_data[140][87] = 11;
        pixel_data[140][88] = 11;
        pixel_data[140][89] = 11;
        pixel_data[140][90] = 11;
        pixel_data[140][91] = 11;
        pixel_data[140][92] = 11;
        pixel_data[140][93] = 11;
        pixel_data[140][94] = 11;
        pixel_data[140][95] = 11;
        pixel_data[140][96] = 11;
        pixel_data[140][97] = 11;
        pixel_data[140][98] = 11;
        pixel_data[140][99] = 11;
        pixel_data[140][100] = 11;
        pixel_data[140][101] = 11;
        pixel_data[140][102] = 11;
        pixel_data[140][103] = 11;
        pixel_data[140][104] = 11;
        pixel_data[140][105] = 11;
        pixel_data[140][106] = 13;
        pixel_data[140][107] = 0;
        pixel_data[140][108] = 0;
        pixel_data[140][109] = 0;
        pixel_data[140][110] = 0;
        pixel_data[140][111] = 0;
        pixel_data[140][112] = 0;
        pixel_data[140][113] = 0;
        pixel_data[140][114] = 0;
        pixel_data[140][115] = 0;
        pixel_data[140][116] = 0;
        pixel_data[140][117] = 0;
        pixel_data[140][118] = 0;
        pixel_data[140][119] = 0;
        pixel_data[140][120] = 0;
        pixel_data[140][121] = 0;
        pixel_data[140][122] = 0;
        pixel_data[140][123] = 0;
        pixel_data[140][124] = 0;
        pixel_data[140][125] = 0;
        pixel_data[140][126] = 0;
        pixel_data[140][127] = 0;
        pixel_data[140][128] = 0;
        pixel_data[140][129] = 0;
        pixel_data[140][130] = 0;
        pixel_data[140][131] = 0;
        pixel_data[140][132] = 0;
        pixel_data[140][133] = 0;
        pixel_data[140][134] = 0;
        pixel_data[140][135] = 0;
        pixel_data[140][136] = 0;
        pixel_data[140][137] = 0;
        pixel_data[140][138] = 0;
        pixel_data[140][139] = 0;
        pixel_data[140][140] = 0;
        pixel_data[140][141] = 0;
        pixel_data[140][142] = 0;
        pixel_data[140][143] = 0;
        pixel_data[140][144] = 0;
        pixel_data[140][145] = 0;
        pixel_data[140][146] = 0;
        pixel_data[140][147] = 0;
        pixel_data[140][148] = 0;
        pixel_data[140][149] = 0;
        pixel_data[140][150] = 0;
        pixel_data[140][151] = 0;
        pixel_data[140][152] = 0;
        pixel_data[140][153] = 0;
        pixel_data[140][154] = 0;
        pixel_data[140][155] = 0;
        pixel_data[140][156] = 0;
        pixel_data[140][157] = 0;
        pixel_data[140][158] = 0;
        pixel_data[140][159] = 0;
        pixel_data[140][160] = 0;
        pixel_data[140][161] = 0;
        pixel_data[140][162] = 0;
        pixel_data[140][163] = 0;
        pixel_data[140][164] = 0;
        pixel_data[140][165] = 0;
        pixel_data[140][166] = 0;
        pixel_data[140][167] = 0;
        pixel_data[140][168] = 0;
        pixel_data[140][169] = 0;
        pixel_data[140][170] = 0;
        pixel_data[140][171] = 0;
        pixel_data[140][172] = 0;
        pixel_data[140][173] = 0;
        pixel_data[140][174] = 0;
        pixel_data[140][175] = 0;
        pixel_data[140][176] = 0;
        pixel_data[140][177] = 0;
        pixel_data[140][178] = 0;
        pixel_data[140][179] = 0;
        pixel_data[140][180] = 0;
        pixel_data[140][181] = 0;
        pixel_data[140][182] = 0;
        pixel_data[140][183] = 0;
        pixel_data[140][184] = 0;
        pixel_data[140][185] = 0;
        pixel_data[140][186] = 0;
        pixel_data[140][187] = 0;
        pixel_data[140][188] = 0;
        pixel_data[140][189] = 0;
        pixel_data[140][190] = 0;
        pixel_data[140][191] = 0;
        pixel_data[140][192] = 0;
        pixel_data[140][193] = 0;
        pixel_data[140][194] = 0;
        pixel_data[140][195] = 0;
        pixel_data[140][196] = 0;
        pixel_data[140][197] = 0;
        pixel_data[140][198] = 0;
        pixel_data[140][199] = 0; // y=140
        pixel_data[141][0] = 0;
        pixel_data[141][1] = 0;
        pixel_data[141][2] = 0;
        pixel_data[141][3] = 0;
        pixel_data[141][4] = 0;
        pixel_data[141][5] = 0;
        pixel_data[141][6] = 0;
        pixel_data[141][7] = 0;
        pixel_data[141][8] = 0;
        pixel_data[141][9] = 0;
        pixel_data[141][10] = 0;
        pixel_data[141][11] = 0;
        pixel_data[141][12] = 0;
        pixel_data[141][13] = 0;
        pixel_data[141][14] = 0;
        pixel_data[141][15] = 0;
        pixel_data[141][16] = 0;
        pixel_data[141][17] = 0;
        pixel_data[141][18] = 0;
        pixel_data[141][19] = 0;
        pixel_data[141][20] = 0;
        pixel_data[141][21] = 0;
        pixel_data[141][22] = 0;
        pixel_data[141][23] = 0;
        pixel_data[141][24] = 0;
        pixel_data[141][25] = 0;
        pixel_data[141][26] = 0;
        pixel_data[141][27] = 0;
        pixel_data[141][28] = 0;
        pixel_data[141][29] = 0;
        pixel_data[141][30] = 0;
        pixel_data[141][31] = 0;
        pixel_data[141][32] = 0;
        pixel_data[141][33] = 0;
        pixel_data[141][34] = 0;
        pixel_data[141][35] = 0;
        pixel_data[141][36] = 0;
        pixel_data[141][37] = 0;
        pixel_data[141][38] = 0;
        pixel_data[141][39] = 0;
        pixel_data[141][40] = 0;
        pixel_data[141][41] = 0;
        pixel_data[141][42] = 0;
        pixel_data[141][43] = 0;
        pixel_data[141][44] = 0;
        pixel_data[141][45] = 0;
        pixel_data[141][46] = 0;
        pixel_data[141][47] = 0;
        pixel_data[141][48] = 0;
        pixel_data[141][49] = 0;
        pixel_data[141][50] = 0;
        pixel_data[141][51] = 0;
        pixel_data[141][52] = 0;
        pixel_data[141][53] = 0;
        pixel_data[141][54] = 0;
        pixel_data[141][55] = 0;
        pixel_data[141][56] = 0;
        pixel_data[141][57] = 0;
        pixel_data[141][58] = 0;
        pixel_data[141][59] = 0;
        pixel_data[141][60] = 0;
        pixel_data[141][61] = 0;
        pixel_data[141][62] = 0;
        pixel_data[141][63] = 0;
        pixel_data[141][64] = 0;
        pixel_data[141][65] = 0;
        pixel_data[141][66] = 0;
        pixel_data[141][67] = 9;
        pixel_data[141][68] = 11;
        pixel_data[141][69] = 11;
        pixel_data[141][70] = 11;
        pixel_data[141][71] = 11;
        pixel_data[141][72] = 9;
        pixel_data[141][73] = 8;
        pixel_data[141][74] = 7;
        pixel_data[141][75] = 6;
        pixel_data[141][76] = 4;
        pixel_data[141][77] = 1;
        pixel_data[141][78] = 1;
        pixel_data[141][79] = 1;
        pixel_data[141][80] = 1;
        pixel_data[141][81] = 1;
        pixel_data[141][82] = 1;
        pixel_data[141][83] = 1;
        pixel_data[141][84] = 1;
        pixel_data[141][85] = 1;
        pixel_data[141][86] = 1;
        pixel_data[141][87] = 1;
        pixel_data[141][88] = 1;
        pixel_data[141][89] = 1;
        pixel_data[141][90] = 1;
        pixel_data[141][91] = 1;
        pixel_data[141][92] = 1;
        pixel_data[141][93] = 1;
        pixel_data[141][94] = 1;
        pixel_data[141][95] = 1;
        pixel_data[141][96] = 1;
        pixel_data[141][97] = 1;
        pixel_data[141][98] = 1;
        pixel_data[141][99] = 1;
        pixel_data[141][100] = 1;
        pixel_data[141][101] = 1;
        pixel_data[141][102] = 1;
        pixel_data[141][103] = 4;
        pixel_data[141][104] = 6;
        pixel_data[141][105] = 7;
        pixel_data[141][106] = 7;
        pixel_data[141][107] = 8;
        pixel_data[141][108] = 8;
        pixel_data[141][109] = 9;
        pixel_data[141][110] = 9;
        pixel_data[141][111] = 11;
        pixel_data[141][112] = 11;
        pixel_data[141][113] = 11;
        pixel_data[141][114] = 11;
        pixel_data[141][115] = 11;
        pixel_data[141][116] = 11;
        pixel_data[141][117] = 11;
        pixel_data[141][118] = 11;
        pixel_data[141][119] = 0;
        pixel_data[141][120] = 0;
        pixel_data[141][121] = 0;
        pixel_data[141][122] = 0;
        pixel_data[141][123] = 0;
        pixel_data[141][124] = 0;
        pixel_data[141][125] = 0;
        pixel_data[141][126] = 0;
        pixel_data[141][127] = 0;
        pixel_data[141][128] = 0;
        pixel_data[141][129] = 0;
        pixel_data[141][130] = 0;
        pixel_data[141][131] = 0;
        pixel_data[141][132] = 0;
        pixel_data[141][133] = 0;
        pixel_data[141][134] = 0;
        pixel_data[141][135] = 0;
        pixel_data[141][136] = 0;
        pixel_data[141][137] = 0;
        pixel_data[141][138] = 0;
        pixel_data[141][139] = 0;
        pixel_data[141][140] = 0;
        pixel_data[141][141] = 0;
        pixel_data[141][142] = 0;
        pixel_data[141][143] = 0;
        pixel_data[141][144] = 0;
        pixel_data[141][145] = 0;
        pixel_data[141][146] = 0;
        pixel_data[141][147] = 0;
        pixel_data[141][148] = 0;
        pixel_data[141][149] = 0;
        pixel_data[141][150] = 0;
        pixel_data[141][151] = 0;
        pixel_data[141][152] = 0;
        pixel_data[141][153] = 0;
        pixel_data[141][154] = 0;
        pixel_data[141][155] = 0;
        pixel_data[141][156] = 0;
        pixel_data[141][157] = 0;
        pixel_data[141][158] = 0;
        pixel_data[141][159] = 0;
        pixel_data[141][160] = 0;
        pixel_data[141][161] = 0;
        pixel_data[141][162] = 0;
        pixel_data[141][163] = 0;
        pixel_data[141][164] = 0;
        pixel_data[141][165] = 0;
        pixel_data[141][166] = 0;
        pixel_data[141][167] = 0;
        pixel_data[141][168] = 0;
        pixel_data[141][169] = 0;
        pixel_data[141][170] = 0;
        pixel_data[141][171] = 0;
        pixel_data[141][172] = 0;
        pixel_data[141][173] = 0;
        pixel_data[141][174] = 0;
        pixel_data[141][175] = 0;
        pixel_data[141][176] = 0;
        pixel_data[141][177] = 0;
        pixel_data[141][178] = 0;
        pixel_data[141][179] = 0;
        pixel_data[141][180] = 0;
        pixel_data[141][181] = 0;
        pixel_data[141][182] = 0;
        pixel_data[141][183] = 0;
        pixel_data[141][184] = 0;
        pixel_data[141][185] = 0;
        pixel_data[141][186] = 0;
        pixel_data[141][187] = 0;
        pixel_data[141][188] = 0;
        pixel_data[141][189] = 0;
        pixel_data[141][190] = 0;
        pixel_data[141][191] = 0;
        pixel_data[141][192] = 0;
        pixel_data[141][193] = 0;
        pixel_data[141][194] = 0;
        pixel_data[141][195] = 0;
        pixel_data[141][196] = 0;
        pixel_data[141][197] = 0;
        pixel_data[141][198] = 0;
        pixel_data[141][199] = 0; // y=141
        pixel_data[142][0] = 0;
        pixel_data[142][1] = 0;
        pixel_data[142][2] = 0;
        pixel_data[142][3] = 0;
        pixel_data[142][4] = 0;
        pixel_data[142][5] = 0;
        pixel_data[142][6] = 0;
        pixel_data[142][7] = 0;
        pixel_data[142][8] = 0;
        pixel_data[142][9] = 0;
        pixel_data[142][10] = 0;
        pixel_data[142][11] = 0;
        pixel_data[142][12] = 0;
        pixel_data[142][13] = 0;
        pixel_data[142][14] = 0;
        pixel_data[142][15] = 0;
        pixel_data[142][16] = 0;
        pixel_data[142][17] = 0;
        pixel_data[142][18] = 0;
        pixel_data[142][19] = 0;
        pixel_data[142][20] = 0;
        pixel_data[142][21] = 0;
        pixel_data[142][22] = 0;
        pixel_data[142][23] = 0;
        pixel_data[142][24] = 0;
        pixel_data[142][25] = 0;
        pixel_data[142][26] = 0;
        pixel_data[142][27] = 0;
        pixel_data[142][28] = 0;
        pixel_data[142][29] = 0;
        pixel_data[142][30] = 0;
        pixel_data[142][31] = 0;
        pixel_data[142][32] = 0;
        pixel_data[142][33] = 0;
        pixel_data[142][34] = 0;
        pixel_data[142][35] = 0;
        pixel_data[142][36] = 0;
        pixel_data[142][37] = 0;
        pixel_data[142][38] = 0;
        pixel_data[142][39] = 0;
        pixel_data[142][40] = 0;
        pixel_data[142][41] = 0;
        pixel_data[142][42] = 0;
        pixel_data[142][43] = 0;
        pixel_data[142][44] = 0;
        pixel_data[142][45] = 0;
        pixel_data[142][46] = 0;
        pixel_data[142][47] = 0;
        pixel_data[142][48] = 0;
        pixel_data[142][49] = 0;
        pixel_data[142][50] = 0;
        pixel_data[142][51] = 0;
        pixel_data[142][52] = 0;
        pixel_data[142][53] = 0;
        pixel_data[142][54] = 0;
        pixel_data[142][55] = 0;
        pixel_data[142][56] = 0;
        pixel_data[142][57] = 0;
        pixel_data[142][58] = 0;
        pixel_data[142][59] = 0;
        pixel_data[142][60] = 10;
        pixel_data[142][61] = 11;
        pixel_data[142][62] = 11;
        pixel_data[142][63] = 11;
        pixel_data[142][64] = 11;
        pixel_data[142][65] = 9;
        pixel_data[142][66] = 8;
        pixel_data[142][67] = 7;
        pixel_data[142][68] = 6;
        pixel_data[142][69] = 5;
        pixel_data[142][70] = 1;
        pixel_data[142][71] = 1;
        pixel_data[142][72] = 1;
        pixel_data[142][73] = 1;
        pixel_data[142][74] = 1;
        pixel_data[142][75] = 2;
        pixel_data[142][76] = 2;
        pixel_data[142][77] = 4;
        pixel_data[142][78] = 4;
        pixel_data[142][79] = 4;
        pixel_data[142][80] = 4;
        pixel_data[142][81] = 2;
        pixel_data[142][82] = 1;
        pixel_data[142][83] = 1;
        pixel_data[142][84] = 1;
        pixel_data[142][85] = 1;
        pixel_data[142][86] = 1;
        pixel_data[142][87] = 1;
        pixel_data[142][88] = 1;
        pixel_data[142][89] = 1;
        pixel_data[142][90] = 1;
        pixel_data[142][91] = 1;
        pixel_data[142][92] = 1;
        pixel_data[142][93] = 1;
        pixel_data[142][94] = 1;
        pixel_data[142][95] = 1;
        pixel_data[142][96] = 1;
        pixel_data[142][97] = 1;
        pixel_data[142][98] = 1;
        pixel_data[142][99] = 1;
        pixel_data[142][100] = 1;
        pixel_data[142][101] = 1;
        pixel_data[142][102] = 1;
        pixel_data[142][103] = 1;
        pixel_data[142][104] = 1;
        pixel_data[142][105] = 1;
        pixel_data[142][106] = 1;
        pixel_data[142][107] = 1;
        pixel_data[142][108] = 1;
        pixel_data[142][109] = 1;
        pixel_data[142][110] = 1;
        pixel_data[142][111] = 1;
        pixel_data[142][112] = 1;
        pixel_data[142][113] = 1;
        pixel_data[142][114] = 1;
        pixel_data[142][115] = 4;
        pixel_data[142][116] = 5;
        pixel_data[142][117] = 7;
        pixel_data[142][118] = 8;
        pixel_data[142][119] = 8;
        pixel_data[142][120] = 9;
        pixel_data[142][121] = 11;
        pixel_data[142][122] = 11;
        pixel_data[142][123] = 11;
        pixel_data[142][124] = 11;
        pixel_data[142][125] = 11;
        pixel_data[142][126] = 11;
        pixel_data[142][127] = 0;
        pixel_data[142][128] = 0;
        pixel_data[142][129] = 0;
        pixel_data[142][130] = 0;
        pixel_data[142][131] = 0;
        pixel_data[142][132] = 0;
        pixel_data[142][133] = 0;
        pixel_data[142][134] = 0;
        pixel_data[142][135] = 0;
        pixel_data[142][136] = 0;
        pixel_data[142][137] = 0;
        pixel_data[142][138] = 0;
        pixel_data[142][139] = 0;
        pixel_data[142][140] = 0;
        pixel_data[142][141] = 0;
        pixel_data[142][142] = 0;
        pixel_data[142][143] = 0;
        pixel_data[142][144] = 0;
        pixel_data[142][145] = 0;
        pixel_data[142][146] = 0;
        pixel_data[142][147] = 0;
        pixel_data[142][148] = 0;
        pixel_data[142][149] = 0;
        pixel_data[142][150] = 0;
        pixel_data[142][151] = 0;
        pixel_data[142][152] = 0;
        pixel_data[142][153] = 0;
        pixel_data[142][154] = 0;
        pixel_data[142][155] = 0;
        pixel_data[142][156] = 0;
        pixel_data[142][157] = 0;
        pixel_data[142][158] = 0;
        pixel_data[142][159] = 0;
        pixel_data[142][160] = 0;
        pixel_data[142][161] = 0;
        pixel_data[142][162] = 0;
        pixel_data[142][163] = 0;
        pixel_data[142][164] = 0;
        pixel_data[142][165] = 0;
        pixel_data[142][166] = 0;
        pixel_data[142][167] = 0;
        pixel_data[142][168] = 0;
        pixel_data[142][169] = 0;
        pixel_data[142][170] = 0;
        pixel_data[142][171] = 0;
        pixel_data[142][172] = 0;
        pixel_data[142][173] = 0;
        pixel_data[142][174] = 0;
        pixel_data[142][175] = 0;
        pixel_data[142][176] = 0;
        pixel_data[142][177] = 0;
        pixel_data[142][178] = 0;
        pixel_data[142][179] = 0;
        pixel_data[142][180] = 0;
        pixel_data[142][181] = 0;
        pixel_data[142][182] = 0;
        pixel_data[142][183] = 0;
        pixel_data[142][184] = 0;
        pixel_data[142][185] = 0;
        pixel_data[142][186] = 0;
        pixel_data[142][187] = 0;
        pixel_data[142][188] = 0;
        pixel_data[142][189] = 0;
        pixel_data[142][190] = 0;
        pixel_data[142][191] = 0;
        pixel_data[142][192] = 0;
        pixel_data[142][193] = 0;
        pixel_data[142][194] = 0;
        pixel_data[142][195] = 0;
        pixel_data[142][196] = 0;
        pixel_data[142][197] = 0;
        pixel_data[142][198] = 0;
        pixel_data[142][199] = 0; // y=142
        pixel_data[143][0] = 0;
        pixel_data[143][1] = 0;
        pixel_data[143][2] = 0;
        pixel_data[143][3] = 0;
        pixel_data[143][4] = 0;
        pixel_data[143][5] = 0;
        pixel_data[143][6] = 0;
        pixel_data[143][7] = 0;
        pixel_data[143][8] = 0;
        pixel_data[143][9] = 0;
        pixel_data[143][10] = 0;
        pixel_data[143][11] = 0;
        pixel_data[143][12] = 0;
        pixel_data[143][13] = 0;
        pixel_data[143][14] = 0;
        pixel_data[143][15] = 0;
        pixel_data[143][16] = 0;
        pixel_data[143][17] = 0;
        pixel_data[143][18] = 0;
        pixel_data[143][19] = 0;
        pixel_data[143][20] = 0;
        pixel_data[143][21] = 0;
        pixel_data[143][22] = 0;
        pixel_data[143][23] = 0;
        pixel_data[143][24] = 0;
        pixel_data[143][25] = 0;
        pixel_data[143][26] = 0;
        pixel_data[143][27] = 0;
        pixel_data[143][28] = 0;
        pixel_data[143][29] = 0;
        pixel_data[143][30] = 0;
        pixel_data[143][31] = 0;
        pixel_data[143][32] = 0;
        pixel_data[143][33] = 0;
        pixel_data[143][34] = 0;
        pixel_data[143][35] = 0;
        pixel_data[143][36] = 0;
        pixel_data[143][37] = 0;
        pixel_data[143][38] = 0;
        pixel_data[143][39] = 0;
        pixel_data[143][40] = 0;
        pixel_data[143][41] = 0;
        pixel_data[143][42] = 0;
        pixel_data[143][43] = 0;
        pixel_data[143][44] = 0;
        pixel_data[143][45] = 0;
        pixel_data[143][46] = 0;
        pixel_data[143][47] = 0;
        pixel_data[143][48] = 0;
        pixel_data[143][49] = 0;
        pixel_data[143][50] = 0;
        pixel_data[143][51] = 0;
        pixel_data[143][52] = 0;
        pixel_data[143][53] = 11;
        pixel_data[143][54] = 11;
        pixel_data[143][55] = 11;
        pixel_data[143][56] = 9;
        pixel_data[143][57] = 9;
        pixel_data[143][58] = 8;
        pixel_data[143][59] = 6;
        pixel_data[143][60] = 4;
        pixel_data[143][61] = 1;
        pixel_data[143][62] = 1;
        pixel_data[143][63] = 1;
        pixel_data[143][64] = 1;
        pixel_data[143][65] = 1;
        pixel_data[143][66] = 2;
        pixel_data[143][67] = 4;
        pixel_data[143][68] = 4;
        pixel_data[143][69] = 4;
        pixel_data[143][70] = 4;
        pixel_data[143][71] = 2;
        pixel_data[143][72] = 1;
        pixel_data[143][73] = 1;
        pixel_data[143][74] = 1;
        pixel_data[143][75] = 1;
        pixel_data[143][76] = 1;
        pixel_data[143][77] = 1;
        pixel_data[143][78] = 1;
        pixel_data[143][79] = 1;
        pixel_data[143][80] = 1;
        pixel_data[143][81] = 1;
        pixel_data[143][82] = 1;
        pixel_data[143][83] = 1;
        pixel_data[143][84] = 1;
        pixel_data[143][85] = 1;
        pixel_data[143][86] = 1;
        pixel_data[143][87] = 1;
        pixel_data[143][88] = 1;
        pixel_data[143][89] = 1;
        pixel_data[143][90] = 1;
        pixel_data[143][91] = 1;
        pixel_data[143][92] = 1;
        pixel_data[143][93] = 1;
        pixel_data[143][94] = 1;
        pixel_data[143][95] = 1;
        pixel_data[143][96] = 1;
        pixel_data[143][97] = 1;
        pixel_data[143][98] = 1;
        pixel_data[143][99] = 1;
        pixel_data[143][100] = 1;
        pixel_data[143][101] = 1;
        pixel_data[143][102] = 1;
        pixel_data[143][103] = 1;
        pixel_data[143][104] = 1;
        pixel_data[143][105] = 1;
        pixel_data[143][106] = 1;
        pixel_data[143][107] = 1;
        pixel_data[143][108] = 1;
        pixel_data[143][109] = 1;
        pixel_data[143][110] = 1;
        pixel_data[143][111] = 1;
        pixel_data[143][112] = 1;
        pixel_data[143][113] = 1;
        pixel_data[143][114] = 1;
        pixel_data[143][115] = 1;
        pixel_data[143][116] = 1;
        pixel_data[143][117] = 1;
        pixel_data[143][118] = 1;
        pixel_data[143][119] = 1;
        pixel_data[143][120] = 1;
        pixel_data[143][121] = 1;
        pixel_data[143][122] = 1;
        pixel_data[143][123] = 1;
        pixel_data[143][124] = 1;
        pixel_data[143][125] = 1;
        pixel_data[143][126] = 5;
        pixel_data[143][127] = 7;
        pixel_data[143][128] = 8;
        pixel_data[143][129] = 9;
        pixel_data[143][130] = 11;
        pixel_data[143][131] = 11;
        pixel_data[143][132] = 11;
        pixel_data[143][133] = 11;
        pixel_data[143][134] = 0;
        pixel_data[143][135] = 0;
        pixel_data[143][136] = 0;
        pixel_data[143][137] = 0;
        pixel_data[143][138] = 0;
        pixel_data[143][139] = 0;
        pixel_data[143][140] = 0;
        pixel_data[143][141] = 0;
        pixel_data[143][142] = 0;
        pixel_data[143][143] = 0;
        pixel_data[143][144] = 0;
        pixel_data[143][145] = 0;
        pixel_data[143][146] = 0;
        pixel_data[143][147] = 0;
        pixel_data[143][148] = 0;
        pixel_data[143][149] = 0;
        pixel_data[143][150] = 0;
        pixel_data[143][151] = 0;
        pixel_data[143][152] = 0;
        pixel_data[143][153] = 0;
        pixel_data[143][154] = 0;
        pixel_data[143][155] = 0;
        pixel_data[143][156] = 0;
        pixel_data[143][157] = 0;
        pixel_data[143][158] = 0;
        pixel_data[143][159] = 0;
        pixel_data[143][160] = 0;
        pixel_data[143][161] = 0;
        pixel_data[143][162] = 0;
        pixel_data[143][163] = 0;
        pixel_data[143][164] = 0;
        pixel_data[143][165] = 0;
        pixel_data[143][166] = 0;
        pixel_data[143][167] = 0;
        pixel_data[143][168] = 0;
        pixel_data[143][169] = 0;
        pixel_data[143][170] = 0;
        pixel_data[143][171] = 0;
        pixel_data[143][172] = 0;
        pixel_data[143][173] = 0;
        pixel_data[143][174] = 0;
        pixel_data[143][175] = 0;
        pixel_data[143][176] = 0;
        pixel_data[143][177] = 0;
        pixel_data[143][178] = 0;
        pixel_data[143][179] = 0;
        pixel_data[143][180] = 0;
        pixel_data[143][181] = 0;
        pixel_data[143][182] = 0;
        pixel_data[143][183] = 0;
        pixel_data[143][184] = 0;
        pixel_data[143][185] = 0;
        pixel_data[143][186] = 0;
        pixel_data[143][187] = 0;
        pixel_data[143][188] = 0;
        pixel_data[143][189] = 0;
        pixel_data[143][190] = 0;
        pixel_data[143][191] = 0;
        pixel_data[143][192] = 0;
        pixel_data[143][193] = 0;
        pixel_data[143][194] = 0;
        pixel_data[143][195] = 0;
        pixel_data[143][196] = 0;
        pixel_data[143][197] = 0;
        pixel_data[143][198] = 0;
        pixel_data[143][199] = 0; // y=143
        pixel_data[144][0] = 0;
        pixel_data[144][1] = 0;
        pixel_data[144][2] = 0;
        pixel_data[144][3] = 0;
        pixel_data[144][4] = 0;
        pixel_data[144][5] = 0;
        pixel_data[144][6] = 0;
        pixel_data[144][7] = 0;
        pixel_data[144][8] = 0;
        pixel_data[144][9] = 0;
        pixel_data[144][10] = 0;
        pixel_data[144][11] = 0;
        pixel_data[144][12] = 0;
        pixel_data[144][13] = 0;
        pixel_data[144][14] = 0;
        pixel_data[144][15] = 0;
        pixel_data[144][16] = 0;
        pixel_data[144][17] = 0;
        pixel_data[144][18] = 0;
        pixel_data[144][19] = 0;
        pixel_data[144][20] = 0;
        pixel_data[144][21] = 0;
        pixel_data[144][22] = 0;
        pixel_data[144][23] = 0;
        pixel_data[144][24] = 0;
        pixel_data[144][25] = 0;
        pixel_data[144][26] = 0;
        pixel_data[144][27] = 0;
        pixel_data[144][28] = 0;
        pixel_data[144][29] = 0;
        pixel_data[144][30] = 0;
        pixel_data[144][31] = 0;
        pixel_data[144][32] = 0;
        pixel_data[144][33] = 0;
        pixel_data[144][34] = 0;
        pixel_data[144][35] = 0;
        pixel_data[144][36] = 0;
        pixel_data[144][37] = 0;
        pixel_data[144][38] = 0;
        pixel_data[144][39] = 0;
        pixel_data[144][40] = 0;
        pixel_data[144][41] = 0;
        pixel_data[144][42] = 0;
        pixel_data[144][43] = 0;
        pixel_data[144][44] = 0;
        pixel_data[144][45] = 0;
        pixel_data[144][46] = 0;
        pixel_data[144][47] = 0;
        pixel_data[144][48] = 0;
        pixel_data[144][49] = 11;
        pixel_data[144][50] = 11;
        pixel_data[144][51] = 11;
        pixel_data[144][52] = 9;
        pixel_data[144][53] = 8;
        pixel_data[144][54] = 6;
        pixel_data[144][55] = 4;
        pixel_data[144][56] = 1;
        pixel_data[144][57] = 1;
        pixel_data[144][58] = 1;
        pixel_data[144][59] = 1;
        pixel_data[144][60] = 2;
        pixel_data[144][61] = 4;
        pixel_data[144][62] = 4;
        pixel_data[144][63] = 4;
        pixel_data[144][64] = 4;
        pixel_data[144][65] = 4;
        pixel_data[144][66] = 2;
        pixel_data[144][67] = 1;
        pixel_data[144][68] = 1;
        pixel_data[144][69] = 1;
        pixel_data[144][70] = 1;
        pixel_data[144][71] = 1;
        pixel_data[144][72] = 1;
        pixel_data[144][73] = 1;
        pixel_data[144][74] = 1;
        pixel_data[144][75] = 1;
        pixel_data[144][76] = 1;
        pixel_data[144][77] = 1;
        pixel_data[144][78] = 1;
        pixel_data[144][79] = 1;
        pixel_data[144][80] = 1;
        pixel_data[144][81] = 1;
        pixel_data[144][82] = 1;
        pixel_data[144][83] = 1;
        pixel_data[144][84] = 1;
        pixel_data[144][85] = 1;
        pixel_data[144][86] = 1;
        pixel_data[144][87] = 1;
        pixel_data[144][88] = 1;
        pixel_data[144][89] = 1;
        pixel_data[144][90] = 1;
        pixel_data[144][91] = 1;
        pixel_data[144][92] = 1;
        pixel_data[144][93] = 1;
        pixel_data[144][94] = 1;
        pixel_data[144][95] = 1;
        pixel_data[144][96] = 1;
        pixel_data[144][97] = 1;
        pixel_data[144][98] = 1;
        pixel_data[144][99] = 1;
        pixel_data[144][100] = 1;
        pixel_data[144][101] = 1;
        pixel_data[144][102] = 1;
        pixel_data[144][103] = 1;
        pixel_data[144][104] = 1;
        pixel_data[144][105] = 1;
        pixel_data[144][106] = 1;
        pixel_data[144][107] = 1;
        pixel_data[144][108] = 1;
        pixel_data[144][109] = 1;
        pixel_data[144][110] = 1;
        pixel_data[144][111] = 1;
        pixel_data[144][112] = 1;
        pixel_data[144][113] = 1;
        pixel_data[144][114] = 1;
        pixel_data[144][115] = 1;
        pixel_data[144][116] = 1;
        pixel_data[144][117] = 1;
        pixel_data[144][118] = 1;
        pixel_data[144][119] = 1;
        pixel_data[144][120] = 1;
        pixel_data[144][121] = 1;
        pixel_data[144][122] = 1;
        pixel_data[144][123] = 1;
        pixel_data[144][124] = 1;
        pixel_data[144][125] = 1;
        pixel_data[144][126] = 1;
        pixel_data[144][127] = 1;
        pixel_data[144][128] = 1;
        pixel_data[144][129] = 1;
        pixel_data[144][130] = 1;
        pixel_data[144][131] = 5;
        pixel_data[144][132] = 7;
        pixel_data[144][133] = 8;
        pixel_data[144][134] = 9;
        pixel_data[144][135] = 11;
        pixel_data[144][136] = 11;
        pixel_data[144][137] = 10;
        pixel_data[144][138] = 0;
        pixel_data[144][139] = 0;
        pixel_data[144][140] = 0;
        pixel_data[144][141] = 0;
        pixel_data[144][142] = 0;
        pixel_data[144][143] = 0;
        pixel_data[144][144] = 0;
        pixel_data[144][145] = 0;
        pixel_data[144][146] = 0;
        pixel_data[144][147] = 0;
        pixel_data[144][148] = 0;
        pixel_data[144][149] = 0;
        pixel_data[144][150] = 0;
        pixel_data[144][151] = 0;
        pixel_data[144][152] = 0;
        pixel_data[144][153] = 0;
        pixel_data[144][154] = 0;
        pixel_data[144][155] = 0;
        pixel_data[144][156] = 0;
        pixel_data[144][157] = 0;
        pixel_data[144][158] = 0;
        pixel_data[144][159] = 0;
        pixel_data[144][160] = 0;
        pixel_data[144][161] = 0;
        pixel_data[144][162] = 0;
        pixel_data[144][163] = 0;
        pixel_data[144][164] = 0;
        pixel_data[144][165] = 0;
        pixel_data[144][166] = 0;
        pixel_data[144][167] = 0;
        pixel_data[144][168] = 0;
        pixel_data[144][169] = 0;
        pixel_data[144][170] = 0;
        pixel_data[144][171] = 0;
        pixel_data[144][172] = 0;
        pixel_data[144][173] = 0;
        pixel_data[144][174] = 0;
        pixel_data[144][175] = 0;
        pixel_data[144][176] = 0;
        pixel_data[144][177] = 0;
        pixel_data[144][178] = 0;
        pixel_data[144][179] = 0;
        pixel_data[144][180] = 0;
        pixel_data[144][181] = 0;
        pixel_data[144][182] = 0;
        pixel_data[144][183] = 0;
        pixel_data[144][184] = 0;
        pixel_data[144][185] = 0;
        pixel_data[144][186] = 0;
        pixel_data[144][187] = 0;
        pixel_data[144][188] = 0;
        pixel_data[144][189] = 0;
        pixel_data[144][190] = 0;
        pixel_data[144][191] = 0;
        pixel_data[144][192] = 0;
        pixel_data[144][193] = 0;
        pixel_data[144][194] = 0;
        pixel_data[144][195] = 0;
        pixel_data[144][196] = 0;
        pixel_data[144][197] = 0;
        pixel_data[144][198] = 0;
        pixel_data[144][199] = 0; // y=144
        pixel_data[145][0] = 0;
        pixel_data[145][1] = 0;
        pixel_data[145][2] = 0;
        pixel_data[145][3] = 0;
        pixel_data[145][4] = 0;
        pixel_data[145][5] = 0;
        pixel_data[145][6] = 0;
        pixel_data[145][7] = 0;
        pixel_data[145][8] = 0;
        pixel_data[145][9] = 0;
        pixel_data[145][10] = 0;
        pixel_data[145][11] = 0;
        pixel_data[145][12] = 0;
        pixel_data[145][13] = 0;
        pixel_data[145][14] = 0;
        pixel_data[145][15] = 0;
        pixel_data[145][16] = 0;
        pixel_data[145][17] = 0;
        pixel_data[145][18] = 0;
        pixel_data[145][19] = 0;
        pixel_data[145][20] = 0;
        pixel_data[145][21] = 0;
        pixel_data[145][22] = 0;
        pixel_data[145][23] = 0;
        pixel_data[145][24] = 0;
        pixel_data[145][25] = 0;
        pixel_data[145][26] = 0;
        pixel_data[145][27] = 0;
        pixel_data[145][28] = 0;
        pixel_data[145][29] = 0;
        pixel_data[145][30] = 0;
        pixel_data[145][31] = 0;
        pixel_data[145][32] = 0;
        pixel_data[145][33] = 0;
        pixel_data[145][34] = 0;
        pixel_data[145][35] = 0;
        pixel_data[145][36] = 0;
        pixel_data[145][37] = 0;
        pixel_data[145][38] = 0;
        pixel_data[145][39] = 0;
        pixel_data[145][40] = 0;
        pixel_data[145][41] = 0;
        pixel_data[145][42] = 0;
        pixel_data[145][43] = 0;
        pixel_data[145][44] = 0;
        pixel_data[145][45] = 13;
        pixel_data[145][46] = 11;
        pixel_data[145][47] = 11;
        pixel_data[145][48] = 9;
        pixel_data[145][49] = 8;
        pixel_data[145][50] = 6;
        pixel_data[145][51] = 4;
        pixel_data[145][52] = 1;
        pixel_data[145][53] = 1;
        pixel_data[145][54] = 1;
        pixel_data[145][55] = 1;
        pixel_data[145][56] = 1;
        pixel_data[145][57] = 1;
        pixel_data[145][58] = 2;
        pixel_data[145][59] = 4;
        pixel_data[145][60] = 2;
        pixel_data[145][61] = 1;
        pixel_data[145][62] = 1;
        pixel_data[145][63] = 1;
        pixel_data[145][64] = 1;
        pixel_data[145][65] = 1;
        pixel_data[145][66] = 1;
        pixel_data[145][67] = 1;
        pixel_data[145][68] = 1;
        pixel_data[145][69] = 1;
        pixel_data[145][70] = 1;
        pixel_data[145][71] = 1;
        pixel_data[145][72] = 1;
        pixel_data[145][73] = 1;
        pixel_data[145][74] = 1;
        pixel_data[145][75] = 1;
        pixel_data[145][76] = 1;
        pixel_data[145][77] = 1;
        pixel_data[145][78] = 1;
        pixel_data[145][79] = 1;
        pixel_data[145][80] = 1;
        pixel_data[145][81] = 1;
        pixel_data[145][82] = 1;
        pixel_data[145][83] = 1;
        pixel_data[145][84] = 1;
        pixel_data[145][85] = 1;
        pixel_data[145][86] = 1;
        pixel_data[145][87] = 1;
        pixel_data[145][88] = 1;
        pixel_data[145][89] = 1;
        pixel_data[145][90] = 1;
        pixel_data[145][91] = 1;
        pixel_data[145][92] = 1;
        pixel_data[145][93] = 1;
        pixel_data[145][94] = 1;
        pixel_data[145][95] = 1;
        pixel_data[145][96] = 1;
        pixel_data[145][97] = 1;
        pixel_data[145][98] = 1;
        pixel_data[145][99] = 1;
        pixel_data[145][100] = 1;
        pixel_data[145][101] = 1;
        pixel_data[145][102] = 1;
        pixel_data[145][103] = 1;
        pixel_data[145][104] = 1;
        pixel_data[145][105] = 1;
        pixel_data[145][106] = 1;
        pixel_data[145][107] = 1;
        pixel_data[145][108] = 1;
        pixel_data[145][109] = 1;
        pixel_data[145][110] = 1;
        pixel_data[145][111] = 1;
        pixel_data[145][112] = 1;
        pixel_data[145][113] = 1;
        pixel_data[145][114] = 1;
        pixel_data[145][115] = 1;
        pixel_data[145][116] = 1;
        pixel_data[145][117] = 1;
        pixel_data[145][118] = 1;
        pixel_data[145][119] = 1;
        pixel_data[145][120] = 1;
        pixel_data[145][121] = 1;
        pixel_data[145][122] = 1;
        pixel_data[145][123] = 1;
        pixel_data[145][124] = 1;
        pixel_data[145][125] = 1;
        pixel_data[145][126] = 1;
        pixel_data[145][127] = 1;
        pixel_data[145][128] = 1;
        pixel_data[145][129] = 1;
        pixel_data[145][130] = 1;
        pixel_data[145][131] = 1;
        pixel_data[145][132] = 1;
        pixel_data[145][133] = 1;
        pixel_data[145][134] = 1;
        pixel_data[145][135] = 4;
        pixel_data[145][136] = 7;
        pixel_data[145][137] = 8;
        pixel_data[145][138] = 9;
        pixel_data[145][139] = 11;
        pixel_data[145][140] = 11;
        pixel_data[145][141] = 13;
        pixel_data[145][142] = 0;
        pixel_data[145][143] = 0;
        pixel_data[145][144] = 0;
        pixel_data[145][145] = 0;
        pixel_data[145][146] = 0;
        pixel_data[145][147] = 0;
        pixel_data[145][148] = 0;
        pixel_data[145][149] = 0;
        pixel_data[145][150] = 0;
        pixel_data[145][151] = 0;
        pixel_data[145][152] = 0;
        pixel_data[145][153] = 0;
        pixel_data[145][154] = 0;
        pixel_data[145][155] = 0;
        pixel_data[145][156] = 0;
        pixel_data[145][157] = 0;
        pixel_data[145][158] = 0;
        pixel_data[145][159] = 0;
        pixel_data[145][160] = 0;
        pixel_data[145][161] = 0;
        pixel_data[145][162] = 0;
        pixel_data[145][163] = 0;
        pixel_data[145][164] = 0;
        pixel_data[145][165] = 0;
        pixel_data[145][166] = 0;
        pixel_data[145][167] = 0;
        pixel_data[145][168] = 0;
        pixel_data[145][169] = 0;
        pixel_data[145][170] = 0;
        pixel_data[145][171] = 0;
        pixel_data[145][172] = 0;
        pixel_data[145][173] = 0;
        pixel_data[145][174] = 0;
        pixel_data[145][175] = 0;
        pixel_data[145][176] = 0;
        pixel_data[145][177] = 0;
        pixel_data[145][178] = 0;
        pixel_data[145][179] = 0;
        pixel_data[145][180] = 0;
        pixel_data[145][181] = 0;
        pixel_data[145][182] = 0;
        pixel_data[145][183] = 0;
        pixel_data[145][184] = 0;
        pixel_data[145][185] = 0;
        pixel_data[145][186] = 0;
        pixel_data[145][187] = 0;
        pixel_data[145][188] = 0;
        pixel_data[145][189] = 0;
        pixel_data[145][190] = 0;
        pixel_data[145][191] = 0;
        pixel_data[145][192] = 0;
        pixel_data[145][193] = 0;
        pixel_data[145][194] = 0;
        pixel_data[145][195] = 0;
        pixel_data[145][196] = 0;
        pixel_data[145][197] = 0;
        pixel_data[145][198] = 0;
        pixel_data[145][199] = 0; // y=145
        pixel_data[146][0] = 0;
        pixel_data[146][1] = 0;
        pixel_data[146][2] = 0;
        pixel_data[146][3] = 0;
        pixel_data[146][4] = 0;
        pixel_data[146][5] = 0;
        pixel_data[146][6] = 0;
        pixel_data[146][7] = 0;
        pixel_data[146][8] = 0;
        pixel_data[146][9] = 0;
        pixel_data[146][10] = 0;
        pixel_data[146][11] = 0;
        pixel_data[146][12] = 0;
        pixel_data[146][13] = 0;
        pixel_data[146][14] = 0;
        pixel_data[146][15] = 0;
        pixel_data[146][16] = 0;
        pixel_data[146][17] = 0;
        pixel_data[146][18] = 0;
        pixel_data[146][19] = 0;
        pixel_data[146][20] = 0;
        pixel_data[146][21] = 0;
        pixel_data[146][22] = 0;
        pixel_data[146][23] = 0;
        pixel_data[146][24] = 0;
        pixel_data[146][25] = 0;
        pixel_data[146][26] = 0;
        pixel_data[146][27] = 0;
        pixel_data[146][28] = 0;
        pixel_data[146][29] = 0;
        pixel_data[146][30] = 0;
        pixel_data[146][31] = 0;
        pixel_data[146][32] = 0;
        pixel_data[146][33] = 0;
        pixel_data[146][34] = 0;
        pixel_data[146][35] = 0;
        pixel_data[146][36] = 0;
        pixel_data[146][37] = 0;
        pixel_data[146][38] = 0;
        pixel_data[146][39] = 0;
        pixel_data[146][40] = 0;
        pixel_data[146][41] = 0;
        pixel_data[146][42] = 11;
        pixel_data[146][43] = 11;
        pixel_data[146][44] = 9;
        pixel_data[146][45] = 8;
        pixel_data[146][46] = 6;
        pixel_data[146][47] = 4;
        pixel_data[146][48] = 4;
        pixel_data[146][49] = 4;
        pixel_data[146][50] = 4;
        pixel_data[146][51] = 4;
        pixel_data[146][52] = 1;
        pixel_data[146][53] = 1;
        pixel_data[146][54] = 1;
        pixel_data[146][55] = 1;
        pixel_data[146][56] = 1;
        pixel_data[146][57] = 1;
        pixel_data[146][58] = 1;
        pixel_data[146][59] = 1;
        pixel_data[146][60] = 1;
        pixel_data[146][61] = 1;
        pixel_data[146][62] = 1;
        pixel_data[146][63] = 1;
        pixel_data[146][64] = 1;
        pixel_data[146][65] = 1;
        pixel_data[146][66] = 1;
        pixel_data[146][67] = 1;
        pixel_data[146][68] = 1;
        pixel_data[146][69] = 1;
        pixel_data[146][70] = 1;
        pixel_data[146][71] = 1;
        pixel_data[146][72] = 1;
        pixel_data[146][73] = 1;
        pixel_data[146][74] = 1;
        pixel_data[146][75] = 1;
        pixel_data[146][76] = 1;
        pixel_data[146][77] = 1;
        pixel_data[146][78] = 1;
        pixel_data[146][79] = 1;
        pixel_data[146][80] = 1;
        pixel_data[146][81] = 1;
        pixel_data[146][82] = 1;
        pixel_data[146][83] = 1;
        pixel_data[146][84] = 1;
        pixel_data[146][85] = 1;
        pixel_data[146][86] = 1;
        pixel_data[146][87] = 1;
        pixel_data[146][88] = 1;
        pixel_data[146][89] = 1;
        pixel_data[146][90] = 1;
        pixel_data[146][91] = 1;
        pixel_data[146][92] = 1;
        pixel_data[146][93] = 1;
        pixel_data[146][94] = 1;
        pixel_data[146][95] = 1;
        pixel_data[146][96] = 1;
        pixel_data[146][97] = 1;
        pixel_data[146][98] = 1;
        pixel_data[146][99] = 1;
        pixel_data[146][100] = 1;
        pixel_data[146][101] = 1;
        pixel_data[146][102] = 1;
        pixel_data[146][103] = 1;
        pixel_data[146][104] = 1;
        pixel_data[146][105] = 1;
        pixel_data[146][106] = 1;
        pixel_data[146][107] = 1;
        pixel_data[146][108] = 1;
        pixel_data[146][109] = 1;
        pixel_data[146][110] = 1;
        pixel_data[146][111] = 1;
        pixel_data[146][112] = 1;
        pixel_data[146][113] = 1;
        pixel_data[146][114] = 1;
        pixel_data[146][115] = 1;
        pixel_data[146][116] = 1;
        pixel_data[146][117] = 1;
        pixel_data[146][118] = 1;
        pixel_data[146][119] = 1;
        pixel_data[146][120] = 1;
        pixel_data[146][121] = 1;
        pixel_data[146][122] = 1;
        pixel_data[146][123] = 1;
        pixel_data[146][124] = 1;
        pixel_data[146][125] = 1;
        pixel_data[146][126] = 1;
        pixel_data[146][127] = 1;
        pixel_data[146][128] = 1;
        pixel_data[146][129] = 1;
        pixel_data[146][130] = 1;
        pixel_data[146][131] = 1;
        pixel_data[146][132] = 1;
        pixel_data[146][133] = 1;
        pixel_data[146][134] = 1;
        pixel_data[146][135] = 1;
        pixel_data[146][136] = 1;
        pixel_data[146][137] = 1;
        pixel_data[146][138] = 1;
        pixel_data[146][139] = 1;
        pixel_data[146][140] = 5;
        pixel_data[146][141] = 7;
        pixel_data[146][142] = 9;
        pixel_data[146][143] = 11;
        pixel_data[146][144] = 11;
        pixel_data[146][145] = 11;
        pixel_data[146][146] = 0;
        pixel_data[146][147] = 0;
        pixel_data[146][148] = 0;
        pixel_data[146][149] = 0;
        pixel_data[146][150] = 0;
        pixel_data[146][151] = 0;
        pixel_data[146][152] = 0;
        pixel_data[146][153] = 0;
        pixel_data[146][154] = 0;
        pixel_data[146][155] = 0;
        pixel_data[146][156] = 0;
        pixel_data[146][157] = 0;
        pixel_data[146][158] = 0;
        pixel_data[146][159] = 0;
        pixel_data[146][160] = 0;
        pixel_data[146][161] = 0;
        pixel_data[146][162] = 0;
        pixel_data[146][163] = 0;
        pixel_data[146][164] = 0;
        pixel_data[146][165] = 0;
        pixel_data[146][166] = 0;
        pixel_data[146][167] = 0;
        pixel_data[146][168] = 0;
        pixel_data[146][169] = 0;
        pixel_data[146][170] = 0;
        pixel_data[146][171] = 0;
        pixel_data[146][172] = 0;
        pixel_data[146][173] = 0;
        pixel_data[146][174] = 0;
        pixel_data[146][175] = 0;
        pixel_data[146][176] = 0;
        pixel_data[146][177] = 0;
        pixel_data[146][178] = 0;
        pixel_data[146][179] = 0;
        pixel_data[146][180] = 0;
        pixel_data[146][181] = 0;
        pixel_data[146][182] = 0;
        pixel_data[146][183] = 0;
        pixel_data[146][184] = 0;
        pixel_data[146][185] = 0;
        pixel_data[146][186] = 0;
        pixel_data[146][187] = 0;
        pixel_data[146][188] = 0;
        pixel_data[146][189] = 0;
        pixel_data[146][190] = 0;
        pixel_data[146][191] = 0;
        pixel_data[146][192] = 0;
        pixel_data[146][193] = 0;
        pixel_data[146][194] = 0;
        pixel_data[146][195] = 0;
        pixel_data[146][196] = 0;
        pixel_data[146][197] = 0;
        pixel_data[146][198] = 0;
        pixel_data[146][199] = 0; // y=146
        pixel_data[147][0] = 0;
        pixel_data[147][1] = 0;
        pixel_data[147][2] = 0;
        pixel_data[147][3] = 0;
        pixel_data[147][4] = 0;
        pixel_data[147][5] = 0;
        pixel_data[147][6] = 0;
        pixel_data[147][7] = 0;
        pixel_data[147][8] = 0;
        pixel_data[147][9] = 0;
        pixel_data[147][10] = 0;
        pixel_data[147][11] = 0;
        pixel_data[147][12] = 0;
        pixel_data[147][13] = 0;
        pixel_data[147][14] = 0;
        pixel_data[147][15] = 0;
        pixel_data[147][16] = 0;
        pixel_data[147][17] = 0;
        pixel_data[147][18] = 0;
        pixel_data[147][19] = 0;
        pixel_data[147][20] = 0;
        pixel_data[147][21] = 0;
        pixel_data[147][22] = 0;
        pixel_data[147][23] = 0;
        pixel_data[147][24] = 0;
        pixel_data[147][25] = 0;
        pixel_data[147][26] = 0;
        pixel_data[147][27] = 0;
        pixel_data[147][28] = 0;
        pixel_data[147][29] = 0;
        pixel_data[147][30] = 0;
        pixel_data[147][31] = 0;
        pixel_data[147][32] = 0;
        pixel_data[147][33] = 0;
        pixel_data[147][34] = 0;
        pixel_data[147][35] = 0;
        pixel_data[147][36] = 0;
        pixel_data[147][37] = 0;
        pixel_data[147][38] = 0;
        pixel_data[147][39] = 0;
        pixel_data[147][40] = 11;
        pixel_data[147][41] = 11;
        pixel_data[147][42] = 9;
        pixel_data[147][43] = 7;
        pixel_data[147][44] = 5;
        pixel_data[147][45] = 4;
        pixel_data[147][46] = 2;
        pixel_data[147][47] = 1;
        pixel_data[147][48] = 1;
        pixel_data[147][49] = 1;
        pixel_data[147][50] = 1;
        pixel_data[147][51] = 1;
        pixel_data[147][52] = 1;
        pixel_data[147][53] = 1;
        pixel_data[147][54] = 1;
        pixel_data[147][55] = 1;
        pixel_data[147][56] = 1;
        pixel_data[147][57] = 1;
        pixel_data[147][58] = 1;
        pixel_data[147][59] = 1;
        pixel_data[147][60] = 1;
        pixel_data[147][61] = 1;
        pixel_data[147][62] = 1;
        pixel_data[147][63] = 1;
        pixel_data[147][64] = 1;
        pixel_data[147][65] = 1;
        pixel_data[147][66] = 1;
        pixel_data[147][67] = 1;
        pixel_data[147][68] = 1;
        pixel_data[147][69] = 1;
        pixel_data[147][70] = 1;
        pixel_data[147][71] = 1;
        pixel_data[147][72] = 1;
        pixel_data[147][73] = 1;
        pixel_data[147][74] = 1;
        pixel_data[147][75] = 1;
        pixel_data[147][76] = 1;
        pixel_data[147][77] = 1;
        pixel_data[147][78] = 1;
        pixel_data[147][79] = 1;
        pixel_data[147][80] = 1;
        pixel_data[147][81] = 1;
        pixel_data[147][82] = 1;
        pixel_data[147][83] = 1;
        pixel_data[147][84] = 1;
        pixel_data[147][85] = 1;
        pixel_data[147][86] = 1;
        pixel_data[147][87] = 1;
        pixel_data[147][88] = 1;
        pixel_data[147][89] = 1;
        pixel_data[147][90] = 1;
        pixel_data[147][91] = 1;
        pixel_data[147][92] = 1;
        pixel_data[147][93] = 1;
        pixel_data[147][94] = 1;
        pixel_data[147][95] = 1;
        pixel_data[147][96] = 1;
        pixel_data[147][97] = 1;
        pixel_data[147][98] = 1;
        pixel_data[147][99] = 1;
        pixel_data[147][100] = 1;
        pixel_data[147][101] = 1;
        pixel_data[147][102] = 1;
        pixel_data[147][103] = 1;
        pixel_data[147][104] = 1;
        pixel_data[147][105] = 1;
        pixel_data[147][106] = 1;
        pixel_data[147][107] = 1;
        pixel_data[147][108] = 1;
        pixel_data[147][109] = 1;
        pixel_data[147][110] = 1;
        pixel_data[147][111] = 1;
        pixel_data[147][112] = 1;
        pixel_data[147][113] = 1;
        pixel_data[147][114] = 1;
        pixel_data[147][115] = 1;
        pixel_data[147][116] = 1;
        pixel_data[147][117] = 1;
        pixel_data[147][118] = 1;
        pixel_data[147][119] = 1;
        pixel_data[147][120] = 1;
        pixel_data[147][121] = 1;
        pixel_data[147][122] = 1;
        pixel_data[147][123] = 1;
        pixel_data[147][124] = 1;
        pixel_data[147][125] = 1;
        pixel_data[147][126] = 1;
        pixel_data[147][127] = 1;
        pixel_data[147][128] = 1;
        pixel_data[147][129] = 1;
        pixel_data[147][130] = 1;
        pixel_data[147][131] = 1;
        pixel_data[147][132] = 1;
        pixel_data[147][133] = 1;
        pixel_data[147][134] = 1;
        pixel_data[147][135] = 1;
        pixel_data[147][136] = 1;
        pixel_data[147][137] = 1;
        pixel_data[147][138] = 1;
        pixel_data[147][139] = 1;
        pixel_data[147][140] = 1;
        pixel_data[147][141] = 1;
        pixel_data[147][142] = 1;
        pixel_data[147][143] = 5;
        pixel_data[147][144] = 7;
        pixel_data[147][145] = 9;
        pixel_data[147][146] = 11;
        pixel_data[147][147] = 11;
        pixel_data[147][148] = 13;
        pixel_data[147][149] = 0;
        pixel_data[147][150] = 0;
        pixel_data[147][151] = 0;
        pixel_data[147][152] = 0;
        pixel_data[147][153] = 0;
        pixel_data[147][154] = 0;
        pixel_data[147][155] = 0;
        pixel_data[147][156] = 0;
        pixel_data[147][157] = 0;
        pixel_data[147][158] = 0;
        pixel_data[147][159] = 0;
        pixel_data[147][160] = 0;
        pixel_data[147][161] = 0;
        pixel_data[147][162] = 0;
        pixel_data[147][163] = 0;
        pixel_data[147][164] = 0;
        pixel_data[147][165] = 0;
        pixel_data[147][166] = 0;
        pixel_data[147][167] = 0;
        pixel_data[147][168] = 0;
        pixel_data[147][169] = 0;
        pixel_data[147][170] = 0;
        pixel_data[147][171] = 0;
        pixel_data[147][172] = 0;
        pixel_data[147][173] = 0;
        pixel_data[147][174] = 0;
        pixel_data[147][175] = 0;
        pixel_data[147][176] = 0;
        pixel_data[147][177] = 0;
        pixel_data[147][178] = 0;
        pixel_data[147][179] = 0;
        pixel_data[147][180] = 0;
        pixel_data[147][181] = 0;
        pixel_data[147][182] = 0;
        pixel_data[147][183] = 0;
        pixel_data[147][184] = 0;
        pixel_data[147][185] = 0;
        pixel_data[147][186] = 0;
        pixel_data[147][187] = 0;
        pixel_data[147][188] = 0;
        pixel_data[147][189] = 0;
        pixel_data[147][190] = 0;
        pixel_data[147][191] = 0;
        pixel_data[147][192] = 0;
        pixel_data[147][193] = 0;
        pixel_data[147][194] = 0;
        pixel_data[147][195] = 0;
        pixel_data[147][196] = 0;
        pixel_data[147][197] = 0;
        pixel_data[147][198] = 0;
        pixel_data[147][199] = 0; // y=147
        pixel_data[148][0] = 0;
        pixel_data[148][1] = 0;
        pixel_data[148][2] = 0;
        pixel_data[148][3] = 0;
        pixel_data[148][4] = 0;
        pixel_data[148][5] = 0;
        pixel_data[148][6] = 0;
        pixel_data[148][7] = 0;
        pixel_data[148][8] = 0;
        pixel_data[148][9] = 0;
        pixel_data[148][10] = 0;
        pixel_data[148][11] = 0;
        pixel_data[148][12] = 0;
        pixel_data[148][13] = 0;
        pixel_data[148][14] = 0;
        pixel_data[148][15] = 0;
        pixel_data[148][16] = 0;
        pixel_data[148][17] = 0;
        pixel_data[148][18] = 0;
        pixel_data[148][19] = 0;
        pixel_data[148][20] = 0;
        pixel_data[148][21] = 0;
        pixel_data[148][22] = 0;
        pixel_data[148][23] = 0;
        pixel_data[148][24] = 0;
        pixel_data[148][25] = 0;
        pixel_data[148][26] = 0;
        pixel_data[148][27] = 0;
        pixel_data[148][28] = 0;
        pixel_data[148][29] = 0;
        pixel_data[148][30] = 0;
        pixel_data[148][31] = 0;
        pixel_data[148][32] = 0;
        pixel_data[148][33] = 0;
        pixel_data[148][34] = 0;
        pixel_data[148][35] = 0;
        pixel_data[148][36] = 0;
        pixel_data[148][37] = 11;
        pixel_data[148][38] = 11;
        pixel_data[148][39] = 9;
        pixel_data[148][40] = 8;
        pixel_data[148][41] = 6;
        pixel_data[148][42] = 1;
        pixel_data[148][43] = 1;
        pixel_data[148][44] = 1;
        pixel_data[148][45] = 1;
        pixel_data[148][46] = 1;
        pixel_data[148][47] = 1;
        pixel_data[148][48] = 1;
        pixel_data[148][49] = 1;
        pixel_data[148][50] = 1;
        pixel_data[148][51] = 1;
        pixel_data[148][52] = 1;
        pixel_data[148][53] = 1;
        pixel_data[148][54] = 1;
        pixel_data[148][55] = 1;
        pixel_data[148][56] = 1;
        pixel_data[148][57] = 1;
        pixel_data[148][58] = 1;
        pixel_data[148][59] = 1;
        pixel_data[148][60] = 1;
        pixel_data[148][61] = 1;
        pixel_data[148][62] = 1;
        pixel_data[148][63] = 1;
        pixel_data[148][64] = 1;
        pixel_data[148][65] = 1;
        pixel_data[148][66] = 1;
        pixel_data[148][67] = 1;
        pixel_data[148][68] = 1;
        pixel_data[148][69] = 1;
        pixel_data[148][70] = 1;
        pixel_data[148][71] = 1;
        pixel_data[148][72] = 1;
        pixel_data[148][73] = 1;
        pixel_data[148][74] = 1;
        pixel_data[148][75] = 1;
        pixel_data[148][76] = 1;
        pixel_data[148][77] = 1;
        pixel_data[148][78] = 1;
        pixel_data[148][79] = 1;
        pixel_data[148][80] = 1;
        pixel_data[148][81] = 1;
        pixel_data[148][82] = 1;
        pixel_data[148][83] = 1;
        pixel_data[148][84] = 1;
        pixel_data[148][85] = 1;
        pixel_data[148][86] = 1;
        pixel_data[148][87] = 1;
        pixel_data[148][88] = 1;
        pixel_data[148][89] = 1;
        pixel_data[148][90] = 1;
        pixel_data[148][91] = 1;
        pixel_data[148][92] = 1;
        pixel_data[148][93] = 1;
        pixel_data[148][94] = 1;
        pixel_data[148][95] = 1;
        pixel_data[148][96] = 1;
        pixel_data[148][97] = 1;
        pixel_data[148][98] = 1;
        pixel_data[148][99] = 1;
        pixel_data[148][100] = 1;
        pixel_data[148][101] = 1;
        pixel_data[148][102] = 1;
        pixel_data[148][103] = 1;
        pixel_data[148][104] = 1;
        pixel_data[148][105] = 1;
        pixel_data[148][106] = 1;
        pixel_data[148][107] = 1;
        pixel_data[148][108] = 1;
        pixel_data[148][109] = 1;
        pixel_data[148][110] = 1;
        pixel_data[148][111] = 1;
        pixel_data[148][112] = 1;
        pixel_data[148][113] = 1;
        pixel_data[148][114] = 1;
        pixel_data[148][115] = 1;
        pixel_data[148][116] = 1;
        pixel_data[148][117] = 1;
        pixel_data[148][118] = 1;
        pixel_data[148][119] = 1;
        pixel_data[148][120] = 1;
        pixel_data[148][121] = 1;
        pixel_data[148][122] = 1;
        pixel_data[148][123] = 1;
        pixel_data[148][124] = 1;
        pixel_data[148][125] = 1;
        pixel_data[148][126] = 1;
        pixel_data[148][127] = 1;
        pixel_data[148][128] = 1;
        pixel_data[148][129] = 1;
        pixel_data[148][130] = 1;
        pixel_data[148][131] = 1;
        pixel_data[148][132] = 1;
        pixel_data[148][133] = 1;
        pixel_data[148][134] = 1;
        pixel_data[148][135] = 1;
        pixel_data[148][136] = 1;
        pixel_data[148][137] = 1;
        pixel_data[148][138] = 1;
        pixel_data[148][139] = 1;
        pixel_data[148][140] = 1;
        pixel_data[148][141] = 1;
        pixel_data[148][142] = 1;
        pixel_data[148][143] = 1;
        pixel_data[148][144] = 1;
        pixel_data[148][145] = 1;
        pixel_data[148][146] = 6;
        pixel_data[148][147] = 8;
        pixel_data[148][148] = 9;
        pixel_data[148][149] = 11;
        pixel_data[148][150] = 11;
        pixel_data[148][151] = 0;
        pixel_data[148][152] = 0;
        pixel_data[148][153] = 0;
        pixel_data[148][154] = 0;
        pixel_data[148][155] = 0;
        pixel_data[148][156] = 0;
        pixel_data[148][157] = 0;
        pixel_data[148][158] = 0;
        pixel_data[148][159] = 0;
        pixel_data[148][160] = 0;
        pixel_data[148][161] = 0;
        pixel_data[148][162] = 0;
        pixel_data[148][163] = 0;
        pixel_data[148][164] = 0;
        pixel_data[148][165] = 0;
        pixel_data[148][166] = 0;
        pixel_data[148][167] = 0;
        pixel_data[148][168] = 0;
        pixel_data[148][169] = 0;
        pixel_data[148][170] = 0;
        pixel_data[148][171] = 0;
        pixel_data[148][172] = 0;
        pixel_data[148][173] = 0;
        pixel_data[148][174] = 0;
        pixel_data[148][175] = 0;
        pixel_data[148][176] = 0;
        pixel_data[148][177] = 0;
        pixel_data[148][178] = 0;
        pixel_data[148][179] = 0;
        pixel_data[148][180] = 0;
        pixel_data[148][181] = 0;
        pixel_data[148][182] = 0;
        pixel_data[148][183] = 0;
        pixel_data[148][184] = 0;
        pixel_data[148][185] = 0;
        pixel_data[148][186] = 0;
        pixel_data[148][187] = 0;
        pixel_data[148][188] = 0;
        pixel_data[148][189] = 0;
        pixel_data[148][190] = 0;
        pixel_data[148][191] = 0;
        pixel_data[148][192] = 0;
        pixel_data[148][193] = 0;
        pixel_data[148][194] = 0;
        pixel_data[148][195] = 0;
        pixel_data[148][196] = 0;
        pixel_data[148][197] = 0;
        pixel_data[148][198] = 0;
        pixel_data[148][199] = 0; // y=148
        pixel_data[149][0] = 0;
        pixel_data[149][1] = 0;
        pixel_data[149][2] = 0;
        pixel_data[149][3] = 0;
        pixel_data[149][4] = 0;
        pixel_data[149][5] = 0;
        pixel_data[149][6] = 0;
        pixel_data[149][7] = 0;
        pixel_data[149][8] = 0;
        pixel_data[149][9] = 0;
        pixel_data[149][10] = 0;
        pixel_data[149][11] = 0;
        pixel_data[149][12] = 0;
        pixel_data[149][13] = 0;
        pixel_data[149][14] = 0;
        pixel_data[149][15] = 0;
        pixel_data[149][16] = 0;
        pixel_data[149][17] = 0;
        pixel_data[149][18] = 0;
        pixel_data[149][19] = 0;
        pixel_data[149][20] = 0;
        pixel_data[149][21] = 0;
        pixel_data[149][22] = 0;
        pixel_data[149][23] = 0;
        pixel_data[149][24] = 0;
        pixel_data[149][25] = 0;
        pixel_data[149][26] = 0;
        pixel_data[149][27] = 0;
        pixel_data[149][28] = 0;
        pixel_data[149][29] = 0;
        pixel_data[149][30] = 0;
        pixel_data[149][31] = 0;
        pixel_data[149][32] = 0;
        pixel_data[149][33] = 0;
        pixel_data[149][34] = 11;
        pixel_data[149][35] = 11;
        pixel_data[149][36] = 11;
        pixel_data[149][37] = 9;
        pixel_data[149][38] = 7;
        pixel_data[149][39] = 5;
        pixel_data[149][40] = 1;
        pixel_data[149][41] = 1;
        pixel_data[149][42] = 1;
        pixel_data[149][43] = 1;
        pixel_data[149][44] = 1;
        pixel_data[149][45] = 1;
        pixel_data[149][46] = 1;
        pixel_data[149][47] = 1;
        pixel_data[149][48] = 1;
        pixel_data[149][49] = 1;
        pixel_data[149][50] = 1;
        pixel_data[149][51] = 1;
        pixel_data[149][52] = 1;
        pixel_data[149][53] = 1;
        pixel_data[149][54] = 1;
        pixel_data[149][55] = 1;
        pixel_data[149][56] = 1;
        pixel_data[149][57] = 1;
        pixel_data[149][58] = 1;
        pixel_data[149][59] = 1;
        pixel_data[149][60] = 1;
        pixel_data[149][61] = 1;
        pixel_data[149][62] = 1;
        pixel_data[149][63] = 1;
        pixel_data[149][64] = 1;
        pixel_data[149][65] = 1;
        pixel_data[149][66] = 1;
        pixel_data[149][67] = 1;
        pixel_data[149][68] = 1;
        pixel_data[149][69] = 1;
        pixel_data[149][70] = 1;
        pixel_data[149][71] = 1;
        pixel_data[149][72] = 1;
        pixel_data[149][73] = 1;
        pixel_data[149][74] = 1;
        pixel_data[149][75] = 1;
        pixel_data[149][76] = 1;
        pixel_data[149][77] = 1;
        pixel_data[149][78] = 1;
        pixel_data[149][79] = 1;
        pixel_data[149][80] = 1;
        pixel_data[149][81] = 1;
        pixel_data[149][82] = 1;
        pixel_data[149][83] = 1;
        pixel_data[149][84] = 1;
        pixel_data[149][85] = 1;
        pixel_data[149][86] = 1;
        pixel_data[149][87] = 1;
        pixel_data[149][88] = 1;
        pixel_data[149][89] = 1;
        pixel_data[149][90] = 1;
        pixel_data[149][91] = 1;
        pixel_data[149][92] = 1;
        pixel_data[149][93] = 1;
        pixel_data[149][94] = 1;
        pixel_data[149][95] = 1;
        pixel_data[149][96] = 1;
        pixel_data[149][97] = 1;
        pixel_data[149][98] = 1;
        pixel_data[149][99] = 1;
        pixel_data[149][100] = 1;
        pixel_data[149][101] = 1;
        pixel_data[149][102] = 1;
        pixel_data[149][103] = 1;
        pixel_data[149][104] = 1;
        pixel_data[149][105] = 1;
        pixel_data[149][106] = 1;
        pixel_data[149][107] = 1;
        pixel_data[149][108] = 1;
        pixel_data[149][109] = 1;
        pixel_data[149][110] = 1;
        pixel_data[149][111] = 1;
        pixel_data[149][112] = 1;
        pixel_data[149][113] = 1;
        pixel_data[149][114] = 1;
        pixel_data[149][115] = 1;
        pixel_data[149][116] = 1;
        pixel_data[149][117] = 1;
        pixel_data[149][118] = 1;
        pixel_data[149][119] = 1;
        pixel_data[149][120] = 1;
        pixel_data[149][121] = 1;
        pixel_data[149][122] = 1;
        pixel_data[149][123] = 1;
        pixel_data[149][124] = 1;
        pixel_data[149][125] = 1;
        pixel_data[149][126] = 1;
        pixel_data[149][127] = 1;
        pixel_data[149][128] = 1;
        pixel_data[149][129] = 1;
        pixel_data[149][130] = 1;
        pixel_data[149][131] = 1;
        pixel_data[149][132] = 1;
        pixel_data[149][133] = 1;
        pixel_data[149][134] = 1;
        pixel_data[149][135] = 1;
        pixel_data[149][136] = 1;
        pixel_data[149][137] = 1;
        pixel_data[149][138] = 1;
        pixel_data[149][139] = 1;
        pixel_data[149][140] = 1;
        pixel_data[149][141] = 1;
        pixel_data[149][142] = 1;
        pixel_data[149][143] = 1;
        pixel_data[149][144] = 1;
        pixel_data[149][145] = 1;
        pixel_data[149][146] = 1;
        pixel_data[149][147] = 1;
        pixel_data[149][148] = 5;
        pixel_data[149][149] = 7;
        pixel_data[149][150] = 9;
        pixel_data[149][151] = 11;
        pixel_data[149][152] = 11;
        pixel_data[149][153] = 13;
        pixel_data[149][154] = 0;
        pixel_data[149][155] = 0;
        pixel_data[149][156] = 0;
        pixel_data[149][157] = 0;
        pixel_data[149][158] = 0;
        pixel_data[149][159] = 0;
        pixel_data[149][160] = 0;
        pixel_data[149][161] = 0;
        pixel_data[149][162] = 0;
        pixel_data[149][163] = 0;
        pixel_data[149][164] = 0;
        pixel_data[149][165] = 0;
        pixel_data[149][166] = 0;
        pixel_data[149][167] = 0;
        pixel_data[149][168] = 0;
        pixel_data[149][169] = 0;
        pixel_data[149][170] = 0;
        pixel_data[149][171] = 0;
        pixel_data[149][172] = 0;
        pixel_data[149][173] = 0;
        pixel_data[149][174] = 0;
        pixel_data[149][175] = 0;
        pixel_data[149][176] = 0;
        pixel_data[149][177] = 0;
        pixel_data[149][178] = 0;
        pixel_data[149][179] = 0;
        pixel_data[149][180] = 0;
        pixel_data[149][181] = 0;
        pixel_data[149][182] = 0;
        pixel_data[149][183] = 0;
        pixel_data[149][184] = 0;
        pixel_data[149][185] = 0;
        pixel_data[149][186] = 0;
        pixel_data[149][187] = 0;
        pixel_data[149][188] = 0;
        pixel_data[149][189] = 0;
        pixel_data[149][190] = 0;
        pixel_data[149][191] = 0;
        pixel_data[149][192] = 0;
        pixel_data[149][193] = 0;
        pixel_data[149][194] = 0;
        pixel_data[149][195] = 0;
        pixel_data[149][196] = 0;
        pixel_data[149][197] = 0;
        pixel_data[149][198] = 0;
        pixel_data[149][199] = 0; // y=149
        pixel_data[150][0] = 0;
        pixel_data[150][1] = 0;
        pixel_data[150][2] = 0;
        pixel_data[150][3] = 0;
        pixel_data[150][4] = 0;
        pixel_data[150][5] = 0;
        pixel_data[150][6] = 0;
        pixel_data[150][7] = 0;
        pixel_data[150][8] = 0;
        pixel_data[150][9] = 0;
        pixel_data[150][10] = 0;
        pixel_data[150][11] = 0;
        pixel_data[150][12] = 0;
        pixel_data[150][13] = 0;
        pixel_data[150][14] = 0;
        pixel_data[150][15] = 0;
        pixel_data[150][16] = 0;
        pixel_data[150][17] = 0;
        pixel_data[150][18] = 0;
        pixel_data[150][19] = 0;
        pixel_data[150][20] = 0;
        pixel_data[150][21] = 0;
        pixel_data[150][22] = 0;
        pixel_data[150][23] = 0;
        pixel_data[150][24] = 0;
        pixel_data[150][25] = 0;
        pixel_data[150][26] = 0;
        pixel_data[150][27] = 0;
        pixel_data[150][28] = 0;
        pixel_data[150][29] = 0;
        pixel_data[150][30] = 13;
        pixel_data[150][31] = 11;
        pixel_data[150][32] = 11;
        pixel_data[150][33] = 11;
        pixel_data[150][34] = 9;
        pixel_data[150][35] = 7;
        pixel_data[150][36] = 5;
        pixel_data[150][37] = 1;
        pixel_data[150][38] = 1;
        pixel_data[150][39] = 1;
        pixel_data[150][40] = 1;
        pixel_data[150][41] = 1;
        pixel_data[150][42] = 1;
        pixel_data[150][43] = 1;
        pixel_data[150][44] = 1;
        pixel_data[150][45] = 1;
        pixel_data[150][46] = 1;
        pixel_data[150][47] = 1;
        pixel_data[150][48] = 1;
        pixel_data[150][49] = 1;
        pixel_data[150][50] = 1;
        pixel_data[150][51] = 1;
        pixel_data[150][52] = 1;
        pixel_data[150][53] = 1;
        pixel_data[150][54] = 1;
        pixel_data[150][55] = 1;
        pixel_data[150][56] = 1;
        pixel_data[150][57] = 1;
        pixel_data[150][58] = 1;
        pixel_data[150][59] = 1;
        pixel_data[150][60] = 1;
        pixel_data[150][61] = 1;
        pixel_data[150][62] = 1;
        pixel_data[150][63] = 1;
        pixel_data[150][64] = 1;
        pixel_data[150][65] = 1;
        pixel_data[150][66] = 1;
        pixel_data[150][67] = 1;
        pixel_data[150][68] = 1;
        pixel_data[150][69] = 1;
        pixel_data[150][70] = 1;
        pixel_data[150][71] = 1;
        pixel_data[150][72] = 1;
        pixel_data[150][73] = 1;
        pixel_data[150][74] = 1;
        pixel_data[150][75] = 1;
        pixel_data[150][76] = 1;
        pixel_data[150][77] = 1;
        pixel_data[150][78] = 1;
        pixel_data[150][79] = 1;
        pixel_data[150][80] = 1;
        pixel_data[150][81] = 1;
        pixel_data[150][82] = 1;
        pixel_data[150][83] = 1;
        pixel_data[150][84] = 1;
        pixel_data[150][85] = 1;
        pixel_data[150][86] = 1;
        pixel_data[150][87] = 1;
        pixel_data[150][88] = 1;
        pixel_data[150][89] = 1;
        pixel_data[150][90] = 1;
        pixel_data[150][91] = 1;
        pixel_data[150][92] = 1;
        pixel_data[150][93] = 1;
        pixel_data[150][94] = 1;
        pixel_data[150][95] = 1;
        pixel_data[150][96] = 1;
        pixel_data[150][97] = 1;
        pixel_data[150][98] = 1;
        pixel_data[150][99] = 1;
        pixel_data[150][100] = 1;
        pixel_data[150][101] = 1;
        pixel_data[150][102] = 1;
        pixel_data[150][103] = 1;
        pixel_data[150][104] = 1;
        pixel_data[150][105] = 1;
        pixel_data[150][106] = 1;
        pixel_data[150][107] = 1;
        pixel_data[150][108] = 1;
        pixel_data[150][109] = 1;
        pixel_data[150][110] = 1;
        pixel_data[150][111] = 1;
        pixel_data[150][112] = 1;
        pixel_data[150][113] = 1;
        pixel_data[150][114] = 1;
        pixel_data[150][115] = 1;
        pixel_data[150][116] = 1;
        pixel_data[150][117] = 1;
        pixel_data[150][118] = 1;
        pixel_data[150][119] = 1;
        pixel_data[150][120] = 1;
        pixel_data[150][121] = 1;
        pixel_data[150][122] = 1;
        pixel_data[150][123] = 1;
        pixel_data[150][124] = 1;
        pixel_data[150][125] = 1;
        pixel_data[150][126] = 1;
        pixel_data[150][127] = 1;
        pixel_data[150][128] = 1;
        pixel_data[150][129] = 1;
        pixel_data[150][130] = 1;
        pixel_data[150][131] = 1;
        pixel_data[150][132] = 1;
        pixel_data[150][133] = 1;
        pixel_data[150][134] = 1;
        pixel_data[150][135] = 1;
        pixel_data[150][136] = 1;
        pixel_data[150][137] = 1;
        pixel_data[150][138] = 1;
        pixel_data[150][139] = 1;
        pixel_data[150][140] = 1;
        pixel_data[150][141] = 1;
        pixel_data[150][142] = 1;
        pixel_data[150][143] = 1;
        pixel_data[150][144] = 1;
        pixel_data[150][145] = 1;
        pixel_data[150][146] = 1;
        pixel_data[150][147] = 1;
        pixel_data[150][148] = 1;
        pixel_data[150][149] = 1;
        pixel_data[150][150] = 1;
        pixel_data[150][151] = 2;
        pixel_data[150][152] = 6;
        pixel_data[150][153] = 8;
        pixel_data[150][154] = 11;
        pixel_data[150][155] = 11;
        pixel_data[150][156] = 11;
        pixel_data[150][157] = 0;
        pixel_data[150][158] = 0;
        pixel_data[150][159] = 0;
        pixel_data[150][160] = 0;
        pixel_data[150][161] = 0;
        pixel_data[150][162] = 0;
        pixel_data[150][163] = 0;
        pixel_data[150][164] = 0;
        pixel_data[150][165] = 0;
        pixel_data[150][166] = 0;
        pixel_data[150][167] = 0;
        pixel_data[150][168] = 0;
        pixel_data[150][169] = 0;
        pixel_data[150][170] = 0;
        pixel_data[150][171] = 0;
        pixel_data[150][172] = 0;
        pixel_data[150][173] = 0;
        pixel_data[150][174] = 0;
        pixel_data[150][175] = 0;
        pixel_data[150][176] = 0;
        pixel_data[150][177] = 0;
        pixel_data[150][178] = 0;
        pixel_data[150][179] = 0;
        pixel_data[150][180] = 0;
        pixel_data[150][181] = 0;
        pixel_data[150][182] = 0;
        pixel_data[150][183] = 0;
        pixel_data[150][184] = 0;
        pixel_data[150][185] = 0;
        pixel_data[150][186] = 0;
        pixel_data[150][187] = 0;
        pixel_data[150][188] = 0;
        pixel_data[150][189] = 0;
        pixel_data[150][190] = 0;
        pixel_data[150][191] = 0;
        pixel_data[150][192] = 0;
        pixel_data[150][193] = 0;
        pixel_data[150][194] = 0;
        pixel_data[150][195] = 0;
        pixel_data[150][196] = 0;
        pixel_data[150][197] = 0;
        pixel_data[150][198] = 0;
        pixel_data[150][199] = 0; // y=150
        pixel_data[151][0] = 0;
        pixel_data[151][1] = 0;
        pixel_data[151][2] = 0;
        pixel_data[151][3] = 0;
        pixel_data[151][4] = 0;
        pixel_data[151][5] = 0;
        pixel_data[151][6] = 0;
        pixel_data[151][7] = 0;
        pixel_data[151][8] = 0;
        pixel_data[151][9] = 0;
        pixel_data[151][10] = 0;
        pixel_data[151][11] = 0;
        pixel_data[151][12] = 0;
        pixel_data[151][13] = 0;
        pixel_data[151][14] = 0;
        pixel_data[151][15] = 0;
        pixel_data[151][16] = 0;
        pixel_data[151][17] = 0;
        pixel_data[151][18] = 0;
        pixel_data[151][19] = 0;
        pixel_data[151][20] = 0;
        pixel_data[151][21] = 0;
        pixel_data[151][22] = 0;
        pixel_data[151][23] = 0;
        pixel_data[151][24] = 0;
        pixel_data[151][25] = 0;
        pixel_data[151][26] = 0;
        pixel_data[151][27] = 0;
        pixel_data[151][28] = 0;
        pixel_data[151][29] = 11;
        pixel_data[151][30] = 11;
        pixel_data[151][31] = 11;
        pixel_data[151][32] = 9;
        pixel_data[151][33] = 7;
        pixel_data[151][34] = 4;
        pixel_data[151][35] = 1;
        pixel_data[151][36] = 1;
        pixel_data[151][37] = 1;
        pixel_data[151][38] = 1;
        pixel_data[151][39] = 1;
        pixel_data[151][40] = 1;
        pixel_data[151][41] = 1;
        pixel_data[151][42] = 1;
        pixel_data[151][43] = 1;
        pixel_data[151][44] = 1;
        pixel_data[151][45] = 1;
        pixel_data[151][46] = 1;
        pixel_data[151][47] = 1;
        pixel_data[151][48] = 1;
        pixel_data[151][49] = 1;
        pixel_data[151][50] = 1;
        pixel_data[151][51] = 1;
        pixel_data[151][52] = 1;
        pixel_data[151][53] = 1;
        pixel_data[151][54] = 1;
        pixel_data[151][55] = 1;
        pixel_data[151][56] = 1;
        pixel_data[151][57] = 1;
        pixel_data[151][58] = 1;
        pixel_data[151][59] = 1;
        pixel_data[151][60] = 1;
        pixel_data[151][61] = 1;
        pixel_data[151][62] = 1;
        pixel_data[151][63] = 1;
        pixel_data[151][64] = 1;
        pixel_data[151][65] = 1;
        pixel_data[151][66] = 1;
        pixel_data[151][67] = 1;
        pixel_data[151][68] = 1;
        pixel_data[151][69] = 1;
        pixel_data[151][70] = 1;
        pixel_data[151][71] = 1;
        pixel_data[151][72] = 1;
        pixel_data[151][73] = 1;
        pixel_data[151][74] = 1;
        pixel_data[151][75] = 1;
        pixel_data[151][76] = 1;
        pixel_data[151][77] = 1;
        pixel_data[151][78] = 1;
        pixel_data[151][79] = 1;
        pixel_data[151][80] = 1;
        pixel_data[151][81] = 1;
        pixel_data[151][82] = 1;
        pixel_data[151][83] = 1;
        pixel_data[151][84] = 1;
        pixel_data[151][85] = 1;
        pixel_data[151][86] = 1;
        pixel_data[151][87] = 1;
        pixel_data[151][88] = 1;
        pixel_data[151][89] = 1;
        pixel_data[151][90] = 1;
        pixel_data[151][91] = 1;
        pixel_data[151][92] = 1;
        pixel_data[151][93] = 1;
        pixel_data[151][94] = 1;
        pixel_data[151][95] = 1;
        pixel_data[151][96] = 1;
        pixel_data[151][97] = 1;
        pixel_data[151][98] = 1;
        pixel_data[151][99] = 1;
        pixel_data[151][100] = 1;
        pixel_data[151][101] = 1;
        pixel_data[151][102] = 1;
        pixel_data[151][103] = 1;
        pixel_data[151][104] = 1;
        pixel_data[151][105] = 1;
        pixel_data[151][106] = 1;
        pixel_data[151][107] = 1;
        pixel_data[151][108] = 1;
        pixel_data[151][109] = 1;
        pixel_data[151][110] = 1;
        pixel_data[151][111] = 1;
        pixel_data[151][112] = 1;
        pixel_data[151][113] = 1;
        pixel_data[151][114] = 1;
        pixel_data[151][115] = 1;
        pixel_data[151][116] = 1;
        pixel_data[151][117] = 1;
        pixel_data[151][118] = 1;
        pixel_data[151][119] = 1;
        pixel_data[151][120] = 1;
        pixel_data[151][121] = 1;
        pixel_data[151][122] = 1;
        pixel_data[151][123] = 1;
        pixel_data[151][124] = 1;
        pixel_data[151][125] = 1;
        pixel_data[151][126] = 1;
        pixel_data[151][127] = 1;
        pixel_data[151][128] = 1;
        pixel_data[151][129] = 1;
        pixel_data[151][130] = 1;
        pixel_data[151][131] = 1;
        pixel_data[151][132] = 1;
        pixel_data[151][133] = 1;
        pixel_data[151][134] = 1;
        pixel_data[151][135] = 1;
        pixel_data[151][136] = 1;
        pixel_data[151][137] = 1;
        pixel_data[151][138] = 1;
        pixel_data[151][139] = 1;
        pixel_data[151][140] = 1;
        pixel_data[151][141] = 1;
        pixel_data[151][142] = 1;
        pixel_data[151][143] = 1;
        pixel_data[151][144] = 1;
        pixel_data[151][145] = 1;
        pixel_data[151][146] = 1;
        pixel_data[151][147] = 1;
        pixel_data[151][148] = 1;
        pixel_data[151][149] = 1;
        pixel_data[151][150] = 1;
        pixel_data[151][151] = 1;
        pixel_data[151][152] = 1;
        pixel_data[151][153] = 1;
        pixel_data[151][154] = 6;
        pixel_data[151][155] = 8;
        pixel_data[151][156] = 9;
        pixel_data[151][157] = 11;
        pixel_data[151][158] = 10;
        pixel_data[151][159] = 0;
        pixel_data[151][160] = 0;
        pixel_data[151][161] = 0;
        pixel_data[151][162] = 0;
        pixel_data[151][163] = 0;
        pixel_data[151][164] = 0;
        pixel_data[151][165] = 0;
        pixel_data[151][166] = 0;
        pixel_data[151][167] = 0;
        pixel_data[151][168] = 0;
        pixel_data[151][169] = 0;
        pixel_data[151][170] = 0;
        pixel_data[151][171] = 0;
        pixel_data[151][172] = 0;
        pixel_data[151][173] = 0;
        pixel_data[151][174] = 0;
        pixel_data[151][175] = 0;
        pixel_data[151][176] = 0;
        pixel_data[151][177] = 0;
        pixel_data[151][178] = 0;
        pixel_data[151][179] = 0;
        pixel_data[151][180] = 0;
        pixel_data[151][181] = 0;
        pixel_data[151][182] = 0;
        pixel_data[151][183] = 0;
        pixel_data[151][184] = 0;
        pixel_data[151][185] = 0;
        pixel_data[151][186] = 0;
        pixel_data[151][187] = 0;
        pixel_data[151][188] = 0;
        pixel_data[151][189] = 0;
        pixel_data[151][190] = 0;
        pixel_data[151][191] = 0;
        pixel_data[151][192] = 0;
        pixel_data[151][193] = 0;
        pixel_data[151][194] = 0;
        pixel_data[151][195] = 0;
        pixel_data[151][196] = 0;
        pixel_data[151][197] = 0;
        pixel_data[151][198] = 0;
        pixel_data[151][199] = 0; // y=151
        pixel_data[152][0] = 0;
        pixel_data[152][1] = 0;
        pixel_data[152][2] = 0;
        pixel_data[152][3] = 0;
        pixel_data[152][4] = 0;
        pixel_data[152][5] = 0;
        pixel_data[152][6] = 0;
        pixel_data[152][7] = 0;
        pixel_data[152][8] = 0;
        pixel_data[152][9] = 0;
        pixel_data[152][10] = 0;
        pixel_data[152][11] = 0;
        pixel_data[152][12] = 0;
        pixel_data[152][13] = 0;
        pixel_data[152][14] = 0;
        pixel_data[152][15] = 0;
        pixel_data[152][16] = 0;
        pixel_data[152][17] = 0;
        pixel_data[152][18] = 0;
        pixel_data[152][19] = 0;
        pixel_data[152][20] = 0;
        pixel_data[152][21] = 0;
        pixel_data[152][22] = 0;
        pixel_data[152][23] = 0;
        pixel_data[152][24] = 0;
        pixel_data[152][25] = 0;
        pixel_data[152][26] = 0;
        pixel_data[152][27] = 11;
        pixel_data[152][28] = 11;
        pixel_data[152][29] = 11;
        pixel_data[152][30] = 9;
        pixel_data[152][31] = 8;
        pixel_data[152][32] = 5;
        pixel_data[152][33] = 1;
        pixel_data[152][34] = 1;
        pixel_data[152][35] = 1;
        pixel_data[152][36] = 1;
        pixel_data[152][37] = 1;
        pixel_data[152][38] = 1;
        pixel_data[152][39] = 1;
        pixel_data[152][40] = 1;
        pixel_data[152][41] = 1;
        pixel_data[152][42] = 1;
        pixel_data[152][43] = 1;
        pixel_data[152][44] = 1;
        pixel_data[152][45] = 1;
        pixel_data[152][46] = 1;
        pixel_data[152][47] = 1;
        pixel_data[152][48] = 1;
        pixel_data[152][49] = 1;
        pixel_data[152][50] = 1;
        pixel_data[152][51] = 1;
        pixel_data[152][52] = 1;
        pixel_data[152][53] = 1;
        pixel_data[152][54] = 1;
        pixel_data[152][55] = 1;
        pixel_data[152][56] = 1;
        pixel_data[152][57] = 1;
        pixel_data[152][58] = 1;
        pixel_data[152][59] = 1;
        pixel_data[152][60] = 1;
        pixel_data[152][61] = 1;
        pixel_data[152][62] = 1;
        pixel_data[152][63] = 1;
        pixel_data[152][64] = 1;
        pixel_data[152][65] = 1;
        pixel_data[152][66] = 1;
        pixel_data[152][67] = 1;
        pixel_data[152][68] = 1;
        pixel_data[152][69] = 1;
        pixel_data[152][70] = 1;
        pixel_data[152][71] = 1;
        pixel_data[152][72] = 1;
        pixel_data[152][73] = 1;
        pixel_data[152][74] = 1;
        pixel_data[152][75] = 1;
        pixel_data[152][76] = 1;
        pixel_data[152][77] = 1;
        pixel_data[152][78] = 1;
        pixel_data[152][79] = 1;
        pixel_data[152][80] = 1;
        pixel_data[152][81] = 1;
        pixel_data[152][82] = 1;
        pixel_data[152][83] = 1;
        pixel_data[152][84] = 1;
        pixel_data[152][85] = 1;
        pixel_data[152][86] = 1;
        pixel_data[152][87] = 1;
        pixel_data[152][88] = 1;
        pixel_data[152][89] = 1;
        pixel_data[152][90] = 1;
        pixel_data[152][91] = 1;
        pixel_data[152][92] = 1;
        pixel_data[152][93] = 1;
        pixel_data[152][94] = 1;
        pixel_data[152][95] = 1;
        pixel_data[152][96] = 1;
        pixel_data[152][97] = 1;
        pixel_data[152][98] = 1;
        pixel_data[152][99] = 1;
        pixel_data[152][100] = 1;
        pixel_data[152][101] = 1;
        pixel_data[152][102] = 1;
        pixel_data[152][103] = 1;
        pixel_data[152][104] = 1;
        pixel_data[152][105] = 1;
        pixel_data[152][106] = 1;
        pixel_data[152][107] = 1;
        pixel_data[152][108] = 1;
        pixel_data[152][109] = 1;
        pixel_data[152][110] = 1;
        pixel_data[152][111] = 1;
        pixel_data[152][112] = 1;
        pixel_data[152][113] = 1;
        pixel_data[152][114] = 1;
        pixel_data[152][115] = 1;
        pixel_data[152][116] = 1;
        pixel_data[152][117] = 1;
        pixel_data[152][118] = 1;
        pixel_data[152][119] = 1;
        pixel_data[152][120] = 1;
        pixel_data[152][121] = 1;
        pixel_data[152][122] = 1;
        pixel_data[152][123] = 1;
        pixel_data[152][124] = 1;
        pixel_data[152][125] = 1;
        pixel_data[152][126] = 1;
        pixel_data[152][127] = 1;
        pixel_data[152][128] = 1;
        pixel_data[152][129] = 1;
        pixel_data[152][130] = 1;
        pixel_data[152][131] = 1;
        pixel_data[152][132] = 1;
        pixel_data[152][133] = 1;
        pixel_data[152][134] = 1;
        pixel_data[152][135] = 1;
        pixel_data[152][136] = 1;
        pixel_data[152][137] = 1;
        pixel_data[152][138] = 1;
        pixel_data[152][139] = 1;
        pixel_data[152][140] = 1;
        pixel_data[152][141] = 1;
        pixel_data[152][142] = 1;
        pixel_data[152][143] = 1;
        pixel_data[152][144] = 1;
        pixel_data[152][145] = 1;
        pixel_data[152][146] = 1;
        pixel_data[152][147] = 1;
        pixel_data[152][148] = 1;
        pixel_data[152][149] = 1;
        pixel_data[152][150] = 1;
        pixel_data[152][151] = 1;
        pixel_data[152][152] = 1;
        pixel_data[152][153] = 1;
        pixel_data[152][154] = 1;
        pixel_data[152][155] = 1;
        pixel_data[152][156] = 5;
        pixel_data[152][157] = 8;
        pixel_data[152][158] = 9;
        pixel_data[152][159] = 11;
        pixel_data[152][160] = 11;
        pixel_data[152][161] = 0;
        pixel_data[152][162] = 0;
        pixel_data[152][163] = 0;
        pixel_data[152][164] = 0;
        pixel_data[152][165] = 0;
        pixel_data[152][166] = 0;
        pixel_data[152][167] = 0;
        pixel_data[152][168] = 0;
        pixel_data[152][169] = 0;
        pixel_data[152][170] = 0;
        pixel_data[152][171] = 0;
        pixel_data[152][172] = 0;
        pixel_data[152][173] = 0;
        pixel_data[152][174] = 0;
        pixel_data[152][175] = 0;
        pixel_data[152][176] = 0;
        pixel_data[152][177] = 0;
        pixel_data[152][178] = 0;
        pixel_data[152][179] = 0;
        pixel_data[152][180] = 0;
        pixel_data[152][181] = 0;
        pixel_data[152][182] = 0;
        pixel_data[152][183] = 0;
        pixel_data[152][184] = 0;
        pixel_data[152][185] = 0;
        pixel_data[152][186] = 0;
        pixel_data[152][187] = 0;
        pixel_data[152][188] = 0;
        pixel_data[152][189] = 0;
        pixel_data[152][190] = 0;
        pixel_data[152][191] = 0;
        pixel_data[152][192] = 0;
        pixel_data[152][193] = 0;
        pixel_data[152][194] = 0;
        pixel_data[152][195] = 0;
        pixel_data[152][196] = 0;
        pixel_data[152][197] = 0;
        pixel_data[152][198] = 0;
        pixel_data[152][199] = 0; // y=152
        pixel_data[153][0] = 0;
        pixel_data[153][1] = 0;
        pixel_data[153][2] = 0;
        pixel_data[153][3] = 0;
        pixel_data[153][4] = 0;
        pixel_data[153][5] = 0;
        pixel_data[153][6] = 0;
        pixel_data[153][7] = 0;
        pixel_data[153][8] = 0;
        pixel_data[153][9] = 0;
        pixel_data[153][10] = 0;
        pixel_data[153][11] = 0;
        pixel_data[153][12] = 0;
        pixel_data[153][13] = 0;
        pixel_data[153][14] = 0;
        pixel_data[153][15] = 0;
        pixel_data[153][16] = 0;
        pixel_data[153][17] = 0;
        pixel_data[153][18] = 0;
        pixel_data[153][19] = 0;
        pixel_data[153][20] = 0;
        pixel_data[153][21] = 0;
        pixel_data[153][22] = 0;
        pixel_data[153][23] = 0;
        pixel_data[153][24] = 0;
        pixel_data[153][25] = 11;
        pixel_data[153][26] = 11;
        pixel_data[153][27] = 11;
        pixel_data[153][28] = 9;
        pixel_data[153][29] = 8;
        pixel_data[153][30] = 5;
        pixel_data[153][31] = 1;
        pixel_data[153][32] = 1;
        pixel_data[153][33] = 1;
        pixel_data[153][34] = 1;
        pixel_data[153][35] = 1;
        pixel_data[153][36] = 1;
        pixel_data[153][37] = 1;
        pixel_data[153][38] = 1;
        pixel_data[153][39] = 1;
        pixel_data[153][40] = 1;
        pixel_data[153][41] = 1;
        pixel_data[153][42] = 1;
        pixel_data[153][43] = 1;
        pixel_data[153][44] = 1;
        pixel_data[153][45] = 1;
        pixel_data[153][46] = 1;
        pixel_data[153][47] = 1;
        pixel_data[153][48] = 1;
        pixel_data[153][49] = 1;
        pixel_data[153][50] = 1;
        pixel_data[153][51] = 1;
        pixel_data[153][52] = 1;
        pixel_data[153][53] = 1;
        pixel_data[153][54] = 1;
        pixel_data[153][55] = 1;
        pixel_data[153][56] = 1;
        pixel_data[153][57] = 1;
        pixel_data[153][58] = 1;
        pixel_data[153][59] = 1;
        pixel_data[153][60] = 1;
        pixel_data[153][61] = 1;
        pixel_data[153][62] = 1;
        pixel_data[153][63] = 1;
        pixel_data[153][64] = 1;
        pixel_data[153][65] = 1;
        pixel_data[153][66] = 1;
        pixel_data[153][67] = 1;
        pixel_data[153][68] = 1;
        pixel_data[153][69] = 1;
        pixel_data[153][70] = 1;
        pixel_data[153][71] = 1;
        pixel_data[153][72] = 1;
        pixel_data[153][73] = 1;
        pixel_data[153][74] = 1;
        pixel_data[153][75] = 1;
        pixel_data[153][76] = 1;
        pixel_data[153][77] = 1;
        pixel_data[153][78] = 1;
        pixel_data[153][79] = 1;
        pixel_data[153][80] = 1;
        pixel_data[153][81] = 1;
        pixel_data[153][82] = 1;
        pixel_data[153][83] = 1;
        pixel_data[153][84] = 1;
        pixel_data[153][85] = 1;
        pixel_data[153][86] = 1;
        pixel_data[153][87] = 1;
        pixel_data[153][88] = 1;
        pixel_data[153][89] = 1;
        pixel_data[153][90] = 1;
        pixel_data[153][91] = 1;
        pixel_data[153][92] = 1;
        pixel_data[153][93] = 1;
        pixel_data[153][94] = 1;
        pixel_data[153][95] = 1;
        pixel_data[153][96] = 1;
        pixel_data[153][97] = 1;
        pixel_data[153][98] = 1;
        pixel_data[153][99] = 1;
        pixel_data[153][100] = 1;
        pixel_data[153][101] = 1;
        pixel_data[153][102] = 1;
        pixel_data[153][103] = 1;
        pixel_data[153][104] = 1;
        pixel_data[153][105] = 1;
        pixel_data[153][106] = 1;
        pixel_data[153][107] = 1;
        pixel_data[153][108] = 1;
        pixel_data[153][109] = 1;
        pixel_data[153][110] = 1;
        pixel_data[153][111] = 1;
        pixel_data[153][112] = 1;
        pixel_data[153][113] = 1;
        pixel_data[153][114] = 1;
        pixel_data[153][115] = 1;
        pixel_data[153][116] = 1;
        pixel_data[153][117] = 1;
        pixel_data[153][118] = 1;
        pixel_data[153][119] = 1;
        pixel_data[153][120] = 1;
        pixel_data[153][121] = 1;
        pixel_data[153][122] = 1;
        pixel_data[153][123] = 1;
        pixel_data[153][124] = 1;
        pixel_data[153][125] = 1;
        pixel_data[153][126] = 1;
        pixel_data[153][127] = 1;
        pixel_data[153][128] = 1;
        pixel_data[153][129] = 1;
        pixel_data[153][130] = 1;
        pixel_data[153][131] = 1;
        pixel_data[153][132] = 1;
        pixel_data[153][133] = 1;
        pixel_data[153][134] = 1;
        pixel_data[153][135] = 1;
        pixel_data[153][136] = 1;
        pixel_data[153][137] = 1;
        pixel_data[153][138] = 1;
        pixel_data[153][139] = 1;
        pixel_data[153][140] = 1;
        pixel_data[153][141] = 1;
        pixel_data[153][142] = 1;
        pixel_data[153][143] = 1;
        pixel_data[153][144] = 1;
        pixel_data[153][145] = 1;
        pixel_data[153][146] = 1;
        pixel_data[153][147] = 1;
        pixel_data[153][148] = 1;
        pixel_data[153][149] = 1;
        pixel_data[153][150] = 1;
        pixel_data[153][151] = 1;
        pixel_data[153][152] = 1;
        pixel_data[153][153] = 1;
        pixel_data[153][154] = 1;
        pixel_data[153][155] = 1;
        pixel_data[153][156] = 1;
        pixel_data[153][157] = 1;
        pixel_data[153][158] = 1;
        pixel_data[153][159] = 7;
        pixel_data[153][160] = 9;
        pixel_data[153][161] = 11;
        pixel_data[153][162] = 11;
        pixel_data[153][163] = 0;
        pixel_data[153][164] = 0;
        pixel_data[153][165] = 0;
        pixel_data[153][166] = 0;
        pixel_data[153][167] = 0;
        pixel_data[153][168] = 0;
        pixel_data[153][169] = 0;
        pixel_data[153][170] = 0;
        pixel_data[153][171] = 0;
        pixel_data[153][172] = 0;
        pixel_data[153][173] = 0;
        pixel_data[153][174] = 0;
        pixel_data[153][175] = 0;
        pixel_data[153][176] = 0;
        pixel_data[153][177] = 0;
        pixel_data[153][178] = 0;
        pixel_data[153][179] = 0;
        pixel_data[153][180] = 0;
        pixel_data[153][181] = 0;
        pixel_data[153][182] = 0;
        pixel_data[153][183] = 0;
        pixel_data[153][184] = 0;
        pixel_data[153][185] = 0;
        pixel_data[153][186] = 0;
        pixel_data[153][187] = 0;
        pixel_data[153][188] = 0;
        pixel_data[153][189] = 0;
        pixel_data[153][190] = 0;
        pixel_data[153][191] = 0;
        pixel_data[153][192] = 0;
        pixel_data[153][193] = 0;
        pixel_data[153][194] = 0;
        pixel_data[153][195] = 0;
        pixel_data[153][196] = 0;
        pixel_data[153][197] = 0;
        pixel_data[153][198] = 0;
        pixel_data[153][199] = 0; // y=153
        pixel_data[154][0] = 0;
        pixel_data[154][1] = 0;
        pixel_data[154][2] = 0;
        pixel_data[154][3] = 0;
        pixel_data[154][4] = 0;
        pixel_data[154][5] = 0;
        pixel_data[154][6] = 0;
        pixel_data[154][7] = 0;
        pixel_data[154][8] = 0;
        pixel_data[154][9] = 0;
        pixel_data[154][10] = 0;
        pixel_data[154][11] = 0;
        pixel_data[154][12] = 0;
        pixel_data[154][13] = 0;
        pixel_data[154][14] = 0;
        pixel_data[154][15] = 0;
        pixel_data[154][16] = 0;
        pixel_data[154][17] = 0;
        pixel_data[154][18] = 0;
        pixel_data[154][19] = 0;
        pixel_data[154][20] = 0;
        pixel_data[154][21] = 0;
        pixel_data[154][22] = 0;
        pixel_data[154][23] = 13;
        pixel_data[154][24] = 11;
        pixel_data[154][25] = 11;
        pixel_data[154][26] = 11;
        pixel_data[154][27] = 8;
        pixel_data[154][28] = 6;
        pixel_data[154][29] = 1;
        pixel_data[154][30] = 1;
        pixel_data[154][31] = 1;
        pixel_data[154][32] = 1;
        pixel_data[154][33] = 1;
        pixel_data[154][34] = 1;
        pixel_data[154][35] = 1;
        pixel_data[154][36] = 1;
        pixel_data[154][37] = 1;
        pixel_data[154][38] = 1;
        pixel_data[154][39] = 1;
        pixel_data[154][40] = 1;
        pixel_data[154][41] = 1;
        pixel_data[154][42] = 1;
        pixel_data[154][43] = 1;
        pixel_data[154][44] = 1;
        pixel_data[154][45] = 1;
        pixel_data[154][46] = 1;
        pixel_data[154][47] = 1;
        pixel_data[154][48] = 1;
        pixel_data[154][49] = 1;
        pixel_data[154][50] = 1;
        pixel_data[154][51] = 1;
        pixel_data[154][52] = 1;
        pixel_data[154][53] = 1;
        pixel_data[154][54] = 1;
        pixel_data[154][55] = 1;
        pixel_data[154][56] = 1;
        pixel_data[154][57] = 1;
        pixel_data[154][58] = 1;
        pixel_data[154][59] = 1;
        pixel_data[154][60] = 1;
        pixel_data[154][61] = 1;
        pixel_data[154][62] = 1;
        pixel_data[154][63] = 1;
        pixel_data[154][64] = 1;
        pixel_data[154][65] = 1;
        pixel_data[154][66] = 1;
        pixel_data[154][67] = 1;
        pixel_data[154][68] = 1;
        pixel_data[154][69] = 1;
        pixel_data[154][70] = 1;
        pixel_data[154][71] = 1;
        pixel_data[154][72] = 1;
        pixel_data[154][73] = 1;
        pixel_data[154][74] = 1;
        pixel_data[154][75] = 1;
        pixel_data[154][76] = 1;
        pixel_data[154][77] = 1;
        pixel_data[154][78] = 1;
        pixel_data[154][79] = 1;
        pixel_data[154][80] = 1;
        pixel_data[154][81] = 1;
        pixel_data[154][82] = 1;
        pixel_data[154][83] = 1;
        pixel_data[154][84] = 1;
        pixel_data[154][85] = 1;
        pixel_data[154][86] = 1;
        pixel_data[154][87] = 1;
        pixel_data[154][88] = 1;
        pixel_data[154][89] = 1;
        pixel_data[154][90] = 1;
        pixel_data[154][91] = 1;
        pixel_data[154][92] = 1;
        pixel_data[154][93] = 1;
        pixel_data[154][94] = 1;
        pixel_data[154][95] = 1;
        pixel_data[154][96] = 1;
        pixel_data[154][97] = 1;
        pixel_data[154][98] = 1;
        pixel_data[154][99] = 1;
        pixel_data[154][100] = 1;
        pixel_data[154][101] = 1;
        pixel_data[154][102] = 1;
        pixel_data[154][103] = 1;
        pixel_data[154][104] = 1;
        pixel_data[154][105] = 1;
        pixel_data[154][106] = 1;
        pixel_data[154][107] = 1;
        pixel_data[154][108] = 1;
        pixel_data[154][109] = 1;
        pixel_data[154][110] = 1;
        pixel_data[154][111] = 1;
        pixel_data[154][112] = 1;
        pixel_data[154][113] = 1;
        pixel_data[154][114] = 1;
        pixel_data[154][115] = 1;
        pixel_data[154][116] = 1;
        pixel_data[154][117] = 1;
        pixel_data[154][118] = 1;
        pixel_data[154][119] = 1;
        pixel_data[154][120] = 1;
        pixel_data[154][121] = 1;
        pixel_data[154][122] = 1;
        pixel_data[154][123] = 1;
        pixel_data[154][124] = 1;
        pixel_data[154][125] = 1;
        pixel_data[154][126] = 1;
        pixel_data[154][127] = 1;
        pixel_data[154][128] = 1;
        pixel_data[154][129] = 1;
        pixel_data[154][130] = 1;
        pixel_data[154][131] = 1;
        pixel_data[154][132] = 1;
        pixel_data[154][133] = 1;
        pixel_data[154][134] = 1;
        pixel_data[154][135] = 1;
        pixel_data[154][136] = 1;
        pixel_data[154][137] = 1;
        pixel_data[154][138] = 1;
        pixel_data[154][139] = 1;
        pixel_data[154][140] = 1;
        pixel_data[154][141] = 1;
        pixel_data[154][142] = 1;
        pixel_data[154][143] = 1;
        pixel_data[154][144] = 1;
        pixel_data[154][145] = 1;
        pixel_data[154][146] = 1;
        pixel_data[154][147] = 1;
        pixel_data[154][148] = 1;
        pixel_data[154][149] = 1;
        pixel_data[154][150] = 1;
        pixel_data[154][151] = 1;
        pixel_data[154][152] = 1;
        pixel_data[154][153] = 1;
        pixel_data[154][154] = 1;
        pixel_data[154][155] = 1;
        pixel_data[154][156] = 1;
        pixel_data[154][157] = 1;
        pixel_data[154][158] = 1;
        pixel_data[154][159] = 1;
        pixel_data[154][160] = 5;
        pixel_data[154][161] = 8;
        pixel_data[154][162] = 9;
        pixel_data[154][163] = 11;
        pixel_data[154][164] = 11;
        pixel_data[154][165] = 0;
        pixel_data[154][166] = 0;
        pixel_data[154][167] = 0;
        pixel_data[154][168] = 0;
        pixel_data[154][169] = 0;
        pixel_data[154][170] = 0;
        pixel_data[154][171] = 0;
        pixel_data[154][172] = 0;
        pixel_data[154][173] = 0;
        pixel_data[154][174] = 0;
        pixel_data[154][175] = 0;
        pixel_data[154][176] = 0;
        pixel_data[154][177] = 0;
        pixel_data[154][178] = 0;
        pixel_data[154][179] = 0;
        pixel_data[154][180] = 0;
        pixel_data[154][181] = 0;
        pixel_data[154][182] = 0;
        pixel_data[154][183] = 0;
        pixel_data[154][184] = 0;
        pixel_data[154][185] = 0;
        pixel_data[154][186] = 0;
        pixel_data[154][187] = 0;
        pixel_data[154][188] = 0;
        pixel_data[154][189] = 0;
        pixel_data[154][190] = 0;
        pixel_data[154][191] = 0;
        pixel_data[154][192] = 0;
        pixel_data[154][193] = 0;
        pixel_data[154][194] = 0;
        pixel_data[154][195] = 0;
        pixel_data[154][196] = 0;
        pixel_data[154][197] = 0;
        pixel_data[154][198] = 0;
        pixel_data[154][199] = 0; // y=154
        pixel_data[155][0] = 0;
        pixel_data[155][1] = 0;
        pixel_data[155][2] = 0;
        pixel_data[155][3] = 0;
        pixel_data[155][4] = 0;
        pixel_data[155][5] = 0;
        pixel_data[155][6] = 0;
        pixel_data[155][7] = 0;
        pixel_data[155][8] = 0;
        pixel_data[155][9] = 0;
        pixel_data[155][10] = 0;
        pixel_data[155][11] = 0;
        pixel_data[155][12] = 0;
        pixel_data[155][13] = 0;
        pixel_data[155][14] = 0;
        pixel_data[155][15] = 0;
        pixel_data[155][16] = 0;
        pixel_data[155][17] = 0;
        pixel_data[155][18] = 0;
        pixel_data[155][19] = 0;
        pixel_data[155][20] = 0;
        pixel_data[155][21] = 0;
        pixel_data[155][22] = 13;
        pixel_data[155][23] = 11;
        pixel_data[155][24] = 11;
        pixel_data[155][25] = 9;
        pixel_data[155][26] = 7;
        pixel_data[155][27] = 2;
        pixel_data[155][28] = 1;
        pixel_data[155][29] = 1;
        pixel_data[155][30] = 1;
        pixel_data[155][31] = 1;
        pixel_data[155][32] = 1;
        pixel_data[155][33] = 1;
        pixel_data[155][34] = 1;
        pixel_data[155][35] = 1;
        pixel_data[155][36] = 1;
        pixel_data[155][37] = 1;
        pixel_data[155][38] = 1;
        pixel_data[155][39] = 1;
        pixel_data[155][40] = 1;
        pixel_data[155][41] = 1;
        pixel_data[155][42] = 1;
        pixel_data[155][43] = 1;
        pixel_data[155][44] = 1;
        pixel_data[155][45] = 1;
        pixel_data[155][46] = 1;
        pixel_data[155][47] = 1;
        pixel_data[155][48] = 1;
        pixel_data[155][49] = 1;
        pixel_data[155][50] = 1;
        pixel_data[155][51] = 1;
        pixel_data[155][52] = 1;
        pixel_data[155][53] = 1;
        pixel_data[155][54] = 1;
        pixel_data[155][55] = 1;
        pixel_data[155][56] = 1;
        pixel_data[155][57] = 1;
        pixel_data[155][58] = 1;
        pixel_data[155][59] = 1;
        pixel_data[155][60] = 1;
        pixel_data[155][61] = 1;
        pixel_data[155][62] = 1;
        pixel_data[155][63] = 1;
        pixel_data[155][64] = 1;
        pixel_data[155][65] = 1;
        pixel_data[155][66] = 1;
        pixel_data[155][67] = 1;
        pixel_data[155][68] = 1;
        pixel_data[155][69] = 1;
        pixel_data[155][70] = 1;
        pixel_data[155][71] = 1;
        pixel_data[155][72] = 1;
        pixel_data[155][73] = 1;
        pixel_data[155][74] = 1;
        pixel_data[155][75] = 1;
        pixel_data[155][76] = 1;
        pixel_data[155][77] = 1;
        pixel_data[155][78] = 1;
        pixel_data[155][79] = 1;
        pixel_data[155][80] = 1;
        pixel_data[155][81] = 1;
        pixel_data[155][82] = 1;
        pixel_data[155][83] = 1;
        pixel_data[155][84] = 1;
        pixel_data[155][85] = 1;
        pixel_data[155][86] = 1;
        pixel_data[155][87] = 1;
        pixel_data[155][88] = 1;
        pixel_data[155][89] = 1;
        pixel_data[155][90] = 1;
        pixel_data[155][91] = 1;
        pixel_data[155][92] = 1;
        pixel_data[155][93] = 1;
        pixel_data[155][94] = 1;
        pixel_data[155][95] = 1;
        pixel_data[155][96] = 1;
        pixel_data[155][97] = 1;
        pixel_data[155][98] = 1;
        pixel_data[155][99] = 1;
        pixel_data[155][100] = 1;
        pixel_data[155][101] = 1;
        pixel_data[155][102] = 1;
        pixel_data[155][103] = 1;
        pixel_data[155][104] = 1;
        pixel_data[155][105] = 1;
        pixel_data[155][106] = 1;
        pixel_data[155][107] = 1;
        pixel_data[155][108] = 1;
        pixel_data[155][109] = 1;
        pixel_data[155][110] = 1;
        pixel_data[155][111] = 1;
        pixel_data[155][112] = 1;
        pixel_data[155][113] = 1;
        pixel_data[155][114] = 1;
        pixel_data[155][115] = 1;
        pixel_data[155][116] = 1;
        pixel_data[155][117] = 1;
        pixel_data[155][118] = 1;
        pixel_data[155][119] = 1;
        pixel_data[155][120] = 1;
        pixel_data[155][121] = 1;
        pixel_data[155][122] = 1;
        pixel_data[155][123] = 1;
        pixel_data[155][124] = 1;
        pixel_data[155][125] = 1;
        pixel_data[155][126] = 1;
        pixel_data[155][127] = 1;
        pixel_data[155][128] = 1;
        pixel_data[155][129] = 1;
        pixel_data[155][130] = 1;
        pixel_data[155][131] = 1;
        pixel_data[155][132] = 1;
        pixel_data[155][133] = 1;
        pixel_data[155][134] = 1;
        pixel_data[155][135] = 1;
        pixel_data[155][136] = 1;
        pixel_data[155][137] = 1;
        pixel_data[155][138] = 1;
        pixel_data[155][139] = 1;
        pixel_data[155][140] = 1;
        pixel_data[155][141] = 1;
        pixel_data[155][142] = 1;
        pixel_data[155][143] = 1;
        pixel_data[155][144] = 1;
        pixel_data[155][145] = 1;
        pixel_data[155][146] = 1;
        pixel_data[155][147] = 1;
        pixel_data[155][148] = 1;
        pixel_data[155][149] = 1;
        pixel_data[155][150] = 1;
        pixel_data[155][151] = 1;
        pixel_data[155][152] = 1;
        pixel_data[155][153] = 1;
        pixel_data[155][154] = 1;
        pixel_data[155][155] = 1;
        pixel_data[155][156] = 1;
        pixel_data[155][157] = 1;
        pixel_data[155][158] = 1;
        pixel_data[155][159] = 1;
        pixel_data[155][160] = 1;
        pixel_data[155][161] = 1;
        pixel_data[155][162] = 6;
        pixel_data[155][163] = 8;
        pixel_data[155][164] = 11;
        pixel_data[155][165] = 11;
        pixel_data[155][166] = 0;
        pixel_data[155][167] = 0;
        pixel_data[155][168] = 0;
        pixel_data[155][169] = 0;
        pixel_data[155][170] = 0;
        pixel_data[155][171] = 0;
        pixel_data[155][172] = 0;
        pixel_data[155][173] = 0;
        pixel_data[155][174] = 0;
        pixel_data[155][175] = 0;
        pixel_data[155][176] = 0;
        pixel_data[155][177] = 0;
        pixel_data[155][178] = 0;
        pixel_data[155][179] = 0;
        pixel_data[155][180] = 0;
        pixel_data[155][181] = 0;
        pixel_data[155][182] = 0;
        pixel_data[155][183] = 0;
        pixel_data[155][184] = 0;
        pixel_data[155][185] = 0;
        pixel_data[155][186] = 0;
        pixel_data[155][187] = 0;
        pixel_data[155][188] = 0;
        pixel_data[155][189] = 0;
        pixel_data[155][190] = 0;
        pixel_data[155][191] = 0;
        pixel_data[155][192] = 0;
        pixel_data[155][193] = 0;
        pixel_data[155][194] = 0;
        pixel_data[155][195] = 0;
        pixel_data[155][196] = 0;
        pixel_data[155][197] = 0;
        pixel_data[155][198] = 0;
        pixel_data[155][199] = 0; // y=155
        pixel_data[156][0] = 0;
        pixel_data[156][1] = 0;
        pixel_data[156][2] = 0;
        pixel_data[156][3] = 0;
        pixel_data[156][4] = 0;
        pixel_data[156][5] = 0;
        pixel_data[156][6] = 0;
        pixel_data[156][7] = 0;
        pixel_data[156][8] = 0;
        pixel_data[156][9] = 0;
        pixel_data[156][10] = 0;
        pixel_data[156][11] = 0;
        pixel_data[156][12] = 0;
        pixel_data[156][13] = 0;
        pixel_data[156][14] = 0;
        pixel_data[156][15] = 0;
        pixel_data[156][16] = 0;
        pixel_data[156][17] = 0;
        pixel_data[156][18] = 0;
        pixel_data[156][19] = 0;
        pixel_data[156][20] = 0;
        pixel_data[156][21] = 11;
        pixel_data[156][22] = 11;
        pixel_data[156][23] = 9;
        pixel_data[156][24] = 7;
        pixel_data[156][25] = 1;
        pixel_data[156][26] = 1;
        pixel_data[156][27] = 1;
        pixel_data[156][28] = 1;
        pixel_data[156][29] = 1;
        pixel_data[156][30] = 1;
        pixel_data[156][31] = 1;
        pixel_data[156][32] = 1;
        pixel_data[156][33] = 1;
        pixel_data[156][34] = 1;
        pixel_data[156][35] = 1;
        pixel_data[156][36] = 1;
        pixel_data[156][37] = 1;
        pixel_data[156][38] = 1;
        pixel_data[156][39] = 1;
        pixel_data[156][40] = 1;
        pixel_data[156][41] = 1;
        pixel_data[156][42] = 1;
        pixel_data[156][43] = 1;
        pixel_data[156][44] = 1;
        pixel_data[156][45] = 1;
        pixel_data[156][46] = 1;
        pixel_data[156][47] = 1;
        pixel_data[156][48] = 1;
        pixel_data[156][49] = 1;
        pixel_data[156][50] = 1;
        pixel_data[156][51] = 1;
        pixel_data[156][52] = 1;
        pixel_data[156][53] = 1;
        pixel_data[156][54] = 1;
        pixel_data[156][55] = 1;
        pixel_data[156][56] = 1;
        pixel_data[156][57] = 1;
        pixel_data[156][58] = 1;
        pixel_data[156][59] = 1;
        pixel_data[156][60] = 1;
        pixel_data[156][61] = 1;
        pixel_data[156][62] = 1;
        pixel_data[156][63] = 1;
        pixel_data[156][64] = 1;
        pixel_data[156][65] = 1;
        pixel_data[156][66] = 1;
        pixel_data[156][67] = 1;
        pixel_data[156][68] = 1;
        pixel_data[156][69] = 1;
        pixel_data[156][70] = 1;
        pixel_data[156][71] = 1;
        pixel_data[156][72] = 1;
        pixel_data[156][73] = 1;
        pixel_data[156][74] = 1;
        pixel_data[156][75] = 1;
        pixel_data[156][76] = 1;
        pixel_data[156][77] = 1;
        pixel_data[156][78] = 1;
        pixel_data[156][79] = 1;
        pixel_data[156][80] = 1;
        pixel_data[156][81] = 1;
        pixel_data[156][82] = 1;
        pixel_data[156][83] = 1;
        pixel_data[156][84] = 1;
        pixel_data[156][85] = 1;
        pixel_data[156][86] = 1;
        pixel_data[156][87] = 1;
        pixel_data[156][88] = 1;
        pixel_data[156][89] = 1;
        pixel_data[156][90] = 1;
        pixel_data[156][91] = 1;
        pixel_data[156][92] = 1;
        pixel_data[156][93] = 1;
        pixel_data[156][94] = 1;
        pixel_data[156][95] = 1;
        pixel_data[156][96] = 1;
        pixel_data[156][97] = 1;
        pixel_data[156][98] = 1;
        pixel_data[156][99] = 1;
        pixel_data[156][100] = 1;
        pixel_data[156][101] = 1;
        pixel_data[156][102] = 1;
        pixel_data[156][103] = 1;
        pixel_data[156][104] = 1;
        pixel_data[156][105] = 1;
        pixel_data[156][106] = 1;
        pixel_data[156][107] = 1;
        pixel_data[156][108] = 1;
        pixel_data[156][109] = 1;
        pixel_data[156][110] = 1;
        pixel_data[156][111] = 1;
        pixel_data[156][112] = 1;
        pixel_data[156][113] = 1;
        pixel_data[156][114] = 1;
        pixel_data[156][115] = 1;
        pixel_data[156][116] = 1;
        pixel_data[156][117] = 1;
        pixel_data[156][118] = 1;
        pixel_data[156][119] = 1;
        pixel_data[156][120] = 1;
        pixel_data[156][121] = 1;
        pixel_data[156][122] = 1;
        pixel_data[156][123] = 1;
        pixel_data[156][124] = 1;
        pixel_data[156][125] = 1;
        pixel_data[156][126] = 1;
        pixel_data[156][127] = 1;
        pixel_data[156][128] = 1;
        pixel_data[156][129] = 1;
        pixel_data[156][130] = 1;
        pixel_data[156][131] = 1;
        pixel_data[156][132] = 1;
        pixel_data[156][133] = 1;
        pixel_data[156][134] = 1;
        pixel_data[156][135] = 1;
        pixel_data[156][136] = 1;
        pixel_data[156][137] = 1;
        pixel_data[156][138] = 1;
        pixel_data[156][139] = 1;
        pixel_data[156][140] = 1;
        pixel_data[156][141] = 1;
        pixel_data[156][142] = 1;
        pixel_data[156][143] = 1;
        pixel_data[156][144] = 1;
        pixel_data[156][145] = 1;
        pixel_data[156][146] = 1;
        pixel_data[156][147] = 1;
        pixel_data[156][148] = 1;
        pixel_data[156][149] = 1;
        pixel_data[156][150] = 1;
        pixel_data[156][151] = 1;
        pixel_data[156][152] = 1;
        pixel_data[156][153] = 1;
        pixel_data[156][154] = 1;
        pixel_data[156][155] = 1;
        pixel_data[156][156] = 1;
        pixel_data[156][157] = 1;
        pixel_data[156][158] = 1;
        pixel_data[156][159] = 1;
        pixel_data[156][160] = 1;
        pixel_data[156][161] = 1;
        pixel_data[156][162] = 1;
        pixel_data[156][163] = 1;
        pixel_data[156][164] = 5;
        pixel_data[156][165] = 8;
        pixel_data[156][166] = 9;
        pixel_data[156][167] = 11;
        pixel_data[156][168] = 11;
        pixel_data[156][169] = 0;
        pixel_data[156][170] = 0;
        pixel_data[156][171] = 0;
        pixel_data[156][172] = 0;
        pixel_data[156][173] = 0;
        pixel_data[156][174] = 0;
        pixel_data[156][175] = 0;
        pixel_data[156][176] = 0;
        pixel_data[156][177] = 0;
        pixel_data[156][178] = 0;
        pixel_data[156][179] = 0;
        pixel_data[156][180] = 0;
        pixel_data[156][181] = 0;
        pixel_data[156][182] = 0;
        pixel_data[156][183] = 0;
        pixel_data[156][184] = 0;
        pixel_data[156][185] = 0;
        pixel_data[156][186] = 0;
        pixel_data[156][187] = 0;
        pixel_data[156][188] = 0;
        pixel_data[156][189] = 0;
        pixel_data[156][190] = 0;
        pixel_data[156][191] = 0;
        pixel_data[156][192] = 0;
        pixel_data[156][193] = 0;
        pixel_data[156][194] = 0;
        pixel_data[156][195] = 0;
        pixel_data[156][196] = 0;
        pixel_data[156][197] = 0;
        pixel_data[156][198] = 0;
        pixel_data[156][199] = 0; // y=156
        pixel_data[157][0] = 0;
        pixel_data[157][1] = 0;
        pixel_data[157][2] = 0;
        pixel_data[157][3] = 0;
        pixel_data[157][4] = 0;
        pixel_data[157][5] = 0;
        pixel_data[157][6] = 0;
        pixel_data[157][7] = 0;
        pixel_data[157][8] = 0;
        pixel_data[157][9] = 0;
        pixel_data[157][10] = 0;
        pixel_data[157][11] = 0;
        pixel_data[157][12] = 0;
        pixel_data[157][13] = 0;
        pixel_data[157][14] = 0;
        pixel_data[157][15] = 0;
        pixel_data[157][16] = 0;
        pixel_data[157][17] = 0;
        pixel_data[157][18] = 0;
        pixel_data[157][19] = 0;
        pixel_data[157][20] = 11;
        pixel_data[157][21] = 11;
        pixel_data[157][22] = 9;
        pixel_data[157][23] = 6;
        pixel_data[157][24] = 1;
        pixel_data[157][25] = 1;
        pixel_data[157][26] = 1;
        pixel_data[157][27] = 1;
        pixel_data[157][28] = 1;
        pixel_data[157][29] = 1;
        pixel_data[157][30] = 1;
        pixel_data[157][31] = 1;
        pixel_data[157][32] = 1;
        pixel_data[157][33] = 1;
        pixel_data[157][34] = 1;
        pixel_data[157][35] = 1;
        pixel_data[157][36] = 1;
        pixel_data[157][37] = 1;
        pixel_data[157][38] = 1;
        pixel_data[157][39] = 1;
        pixel_data[157][40] = 1;
        pixel_data[157][41] = 1;
        pixel_data[157][42] = 1;
        pixel_data[157][43] = 1;
        pixel_data[157][44] = 1;
        pixel_data[157][45] = 1;
        pixel_data[157][46] = 1;
        pixel_data[157][47] = 1;
        pixel_data[157][48] = 1;
        pixel_data[157][49] = 1;
        pixel_data[157][50] = 1;
        pixel_data[157][51] = 1;
        pixel_data[157][52] = 1;
        pixel_data[157][53] = 1;
        pixel_data[157][54] = 1;
        pixel_data[157][55] = 1;
        pixel_data[157][56] = 1;
        pixel_data[157][57] = 1;
        pixel_data[157][58] = 1;
        pixel_data[157][59] = 1;
        pixel_data[157][60] = 1;
        pixel_data[157][61] = 1;
        pixel_data[157][62] = 1;
        pixel_data[157][63] = 1;
        pixel_data[157][64] = 1;
        pixel_data[157][65] = 1;
        pixel_data[157][66] = 1;
        pixel_data[157][67] = 1;
        pixel_data[157][68] = 1;
        pixel_data[157][69] = 1;
        pixel_data[157][70] = 1;
        pixel_data[157][71] = 1;
        pixel_data[157][72] = 1;
        pixel_data[157][73] = 1;
        pixel_data[157][74] = 1;
        pixel_data[157][75] = 1;
        pixel_data[157][76] = 1;
        pixel_data[157][77] = 1;
        pixel_data[157][78] = 1;
        pixel_data[157][79] = 1;
        pixel_data[157][80] = 1;
        pixel_data[157][81] = 1;
        pixel_data[157][82] = 1;
        pixel_data[157][83] = 1;
        pixel_data[157][84] = 1;
        pixel_data[157][85] = 1;
        pixel_data[157][86] = 1;
        pixel_data[157][87] = 1;
        pixel_data[157][88] = 1;
        pixel_data[157][89] = 1;
        pixel_data[157][90] = 1;
        pixel_data[157][91] = 1;
        pixel_data[157][92] = 1;
        pixel_data[157][93] = 1;
        pixel_data[157][94] = 1;
        pixel_data[157][95] = 1;
        pixel_data[157][96] = 1;
        pixel_data[157][97] = 1;
        pixel_data[157][98] = 1;
        pixel_data[157][99] = 1;
        pixel_data[157][100] = 1;
        pixel_data[157][101] = 1;
        pixel_data[157][102] = 1;
        pixel_data[157][103] = 1;
        pixel_data[157][104] = 1;
        pixel_data[157][105] = 1;
        pixel_data[157][106] = 1;
        pixel_data[157][107] = 1;
        pixel_data[157][108] = 1;
        pixel_data[157][109] = 1;
        pixel_data[157][110] = 1;
        pixel_data[157][111] = 1;
        pixel_data[157][112] = 1;
        pixel_data[157][113] = 1;
        pixel_data[157][114] = 1;
        pixel_data[157][115] = 1;
        pixel_data[157][116] = 1;
        pixel_data[157][117] = 1;
        pixel_data[157][118] = 1;
        pixel_data[157][119] = 1;
        pixel_data[157][120] = 1;
        pixel_data[157][121] = 1;
        pixel_data[157][122] = 1;
        pixel_data[157][123] = 1;
        pixel_data[157][124] = 1;
        pixel_data[157][125] = 1;
        pixel_data[157][126] = 1;
        pixel_data[157][127] = 1;
        pixel_data[157][128] = 1;
        pixel_data[157][129] = 1;
        pixel_data[157][130] = 1;
        pixel_data[157][131] = 1;
        pixel_data[157][132] = 1;
        pixel_data[157][133] = 1;
        pixel_data[157][134] = 1;
        pixel_data[157][135] = 1;
        pixel_data[157][136] = 1;
        pixel_data[157][137] = 1;
        pixel_data[157][138] = 1;
        pixel_data[157][139] = 1;
        pixel_data[157][140] = 1;
        pixel_data[157][141] = 1;
        pixel_data[157][142] = 1;
        pixel_data[157][143] = 1;
        pixel_data[157][144] = 1;
        pixel_data[157][145] = 1;
        pixel_data[157][146] = 1;
        pixel_data[157][147] = 1;
        pixel_data[157][148] = 1;
        pixel_data[157][149] = 1;
        pixel_data[157][150] = 1;
        pixel_data[157][151] = 1;
        pixel_data[157][152] = 1;
        pixel_data[157][153] = 1;
        pixel_data[157][154] = 1;
        pixel_data[157][155] = 1;
        pixel_data[157][156] = 1;
        pixel_data[157][157] = 1;
        pixel_data[157][158] = 1;
        pixel_data[157][159] = 1;
        pixel_data[157][160] = 1;
        pixel_data[157][161] = 1;
        pixel_data[157][162] = 1;
        pixel_data[157][163] = 1;
        pixel_data[157][164] = 1;
        pixel_data[157][165] = 1;
        pixel_data[157][166] = 6;
        pixel_data[157][167] = 8;
        pixel_data[157][168] = 11;
        pixel_data[157][169] = 11;
        pixel_data[157][170] = 13;
        pixel_data[157][171] = 0;
        pixel_data[157][172] = 0;
        pixel_data[157][173] = 0;
        pixel_data[157][174] = 0;
        pixel_data[157][175] = 0;
        pixel_data[157][176] = 0;
        pixel_data[157][177] = 0;
        pixel_data[157][178] = 0;
        pixel_data[157][179] = 0;
        pixel_data[157][180] = 0;
        pixel_data[157][181] = 0;
        pixel_data[157][182] = 0;
        pixel_data[157][183] = 0;
        pixel_data[157][184] = 0;
        pixel_data[157][185] = 0;
        pixel_data[157][186] = 0;
        pixel_data[157][187] = 0;
        pixel_data[157][188] = 0;
        pixel_data[157][189] = 0;
        pixel_data[157][190] = 0;
        pixel_data[157][191] = 0;
        pixel_data[157][192] = 0;
        pixel_data[157][193] = 0;
        pixel_data[157][194] = 0;
        pixel_data[157][195] = 0;
        pixel_data[157][196] = 0;
        pixel_data[157][197] = 0;
        pixel_data[157][198] = 0;
        pixel_data[157][199] = 0; // y=157
        pixel_data[158][0] = 0;
        pixel_data[158][1] = 0;
        pixel_data[158][2] = 0;
        pixel_data[158][3] = 0;
        pixel_data[158][4] = 0;
        pixel_data[158][5] = 0;
        pixel_data[158][6] = 0;
        pixel_data[158][7] = 0;
        pixel_data[158][8] = 0;
        pixel_data[158][9] = 0;
        pixel_data[158][10] = 0;
        pixel_data[158][11] = 0;
        pixel_data[158][12] = 0;
        pixel_data[158][13] = 0;
        pixel_data[158][14] = 0;
        pixel_data[158][15] = 0;
        pixel_data[158][16] = 0;
        pixel_data[158][17] = 0;
        pixel_data[158][18] = 0;
        pixel_data[158][19] = 11;
        pixel_data[158][20] = 11;
        pixel_data[158][21] = 8;
        pixel_data[158][22] = 5;
        pixel_data[158][23] = 1;
        pixel_data[158][24] = 1;
        pixel_data[158][25] = 1;
        pixel_data[158][26] = 1;
        pixel_data[158][27] = 1;
        pixel_data[158][28] = 1;
        pixel_data[158][29] = 1;
        pixel_data[158][30] = 1;
        pixel_data[158][31] = 1;
        pixel_data[158][32] = 1;
        pixel_data[158][33] = 1;
        pixel_data[158][34] = 1;
        pixel_data[158][35] = 1;
        pixel_data[158][36] = 1;
        pixel_data[158][37] = 1;
        pixel_data[158][38] = 1;
        pixel_data[158][39] = 1;
        pixel_data[158][40] = 1;
        pixel_data[158][41] = 1;
        pixel_data[158][42] = 1;
        pixel_data[158][43] = 1;
        pixel_data[158][44] = 1;
        pixel_data[158][45] = 1;
        pixel_data[158][46] = 1;
        pixel_data[158][47] = 1;
        pixel_data[158][48] = 1;
        pixel_data[158][49] = 1;
        pixel_data[158][50] = 1;
        pixel_data[158][51] = 1;
        pixel_data[158][52] = 1;
        pixel_data[158][53] = 1;
        pixel_data[158][54] = 1;
        pixel_data[158][55] = 1;
        pixel_data[158][56] = 1;
        pixel_data[158][57] = 1;
        pixel_data[158][58] = 1;
        pixel_data[158][59] = 1;
        pixel_data[158][60] = 1;
        pixel_data[158][61] = 1;
        pixel_data[158][62] = 1;
        pixel_data[158][63] = 1;
        pixel_data[158][64] = 1;
        pixel_data[158][65] = 1;
        pixel_data[158][66] = 1;
        pixel_data[158][67] = 1;
        pixel_data[158][68] = 1;
        pixel_data[158][69] = 1;
        pixel_data[158][70] = 1;
        pixel_data[158][71] = 1;
        pixel_data[158][72] = 1;
        pixel_data[158][73] = 1;
        pixel_data[158][74] = 1;
        pixel_data[158][75] = 1;
        pixel_data[158][76] = 1;
        pixel_data[158][77] = 1;
        pixel_data[158][78] = 1;
        pixel_data[158][79] = 1;
        pixel_data[158][80] = 1;
        pixel_data[158][81] = 1;
        pixel_data[158][82] = 1;
        pixel_data[158][83] = 1;
        pixel_data[158][84] = 1;
        pixel_data[158][85] = 1;
        pixel_data[158][86] = 1;
        pixel_data[158][87] = 1;
        pixel_data[158][88] = 1;
        pixel_data[158][89] = 1;
        pixel_data[158][90] = 1;
        pixel_data[158][91] = 1;
        pixel_data[158][92] = 1;
        pixel_data[158][93] = 1;
        pixel_data[158][94] = 1;
        pixel_data[158][95] = 1;
        pixel_data[158][96] = 1;
        pixel_data[158][97] = 1;
        pixel_data[158][98] = 1;
        pixel_data[158][99] = 1;
        pixel_data[158][100] = 1;
        pixel_data[158][101] = 1;
        pixel_data[158][102] = 1;
        pixel_data[158][103] = 1;
        pixel_data[158][104] = 1;
        pixel_data[158][105] = 1;
        pixel_data[158][106] = 1;
        pixel_data[158][107] = 1;
        pixel_data[158][108] = 1;
        pixel_data[158][109] = 1;
        pixel_data[158][110] = 1;
        pixel_data[158][111] = 1;
        pixel_data[158][112] = 1;
        pixel_data[158][113] = 1;
        pixel_data[158][114] = 1;
        pixel_data[158][115] = 1;
        pixel_data[158][116] = 1;
        pixel_data[158][117] = 1;
        pixel_data[158][118] = 1;
        pixel_data[158][119] = 1;
        pixel_data[158][120] = 1;
        pixel_data[158][121] = 1;
        pixel_data[158][122] = 1;
        pixel_data[158][123] = 1;
        pixel_data[158][124] = 1;
        pixel_data[158][125] = 1;
        pixel_data[158][126] = 1;
        pixel_data[158][127] = 1;
        pixel_data[158][128] = 1;
        pixel_data[158][129] = 1;
        pixel_data[158][130] = 1;
        pixel_data[158][131] = 1;
        pixel_data[158][132] = 1;
        pixel_data[158][133] = 1;
        pixel_data[158][134] = 1;
        pixel_data[158][135] = 1;
        pixel_data[158][136] = 1;
        pixel_data[158][137] = 1;
        pixel_data[158][138] = 1;
        pixel_data[158][139] = 1;
        pixel_data[158][140] = 1;
        pixel_data[158][141] = 1;
        pixel_data[158][142] = 1;
        pixel_data[158][143] = 1;
        pixel_data[158][144] = 1;
        pixel_data[158][145] = 1;
        pixel_data[158][146] = 1;
        pixel_data[158][147] = 1;
        pixel_data[158][148] = 1;
        pixel_data[158][149] = 1;
        pixel_data[158][150] = 1;
        pixel_data[158][151] = 1;
        pixel_data[158][152] = 1;
        pixel_data[158][153] = 1;
        pixel_data[158][154] = 1;
        pixel_data[158][155] = 1;
        pixel_data[158][156] = 1;
        pixel_data[158][157] = 1;
        pixel_data[158][158] = 1;
        pixel_data[158][159] = 1;
        pixel_data[158][160] = 1;
        pixel_data[158][161] = 1;
        pixel_data[158][162] = 1;
        pixel_data[158][163] = 1;
        pixel_data[158][164] = 1;
        pixel_data[158][165] = 1;
        pixel_data[158][166] = 1;
        pixel_data[158][167] = 1;
        pixel_data[158][168] = 7;
        pixel_data[158][169] = 9;
        pixel_data[158][170] = 11;
        pixel_data[158][171] = 11;
        pixel_data[158][172] = 0;
        pixel_data[158][173] = 0;
        pixel_data[158][174] = 0;
        pixel_data[158][175] = 0;
        pixel_data[158][176] = 0;
        pixel_data[158][177] = 0;
        pixel_data[158][178] = 0;
        pixel_data[158][179] = 0;
        pixel_data[158][180] = 0;
        pixel_data[158][181] = 0;
        pixel_data[158][182] = 0;
        pixel_data[158][183] = 0;
        pixel_data[158][184] = 0;
        pixel_data[158][185] = 0;
        pixel_data[158][186] = 0;
        pixel_data[158][187] = 0;
        pixel_data[158][188] = 0;
        pixel_data[158][189] = 0;
        pixel_data[158][190] = 0;
        pixel_data[158][191] = 0;
        pixel_data[158][192] = 0;
        pixel_data[158][193] = 0;
        pixel_data[158][194] = 0;
        pixel_data[158][195] = 0;
        pixel_data[158][196] = 0;
        pixel_data[158][197] = 0;
        pixel_data[158][198] = 0;
        pixel_data[158][199] = 0; // y=158
        pixel_data[159][0] = 0;
        pixel_data[159][1] = 0;
        pixel_data[159][2] = 0;
        pixel_data[159][3] = 0;
        pixel_data[159][4] = 0;
        pixel_data[159][5] = 0;
        pixel_data[159][6] = 0;
        pixel_data[159][7] = 0;
        pixel_data[159][8] = 0;
        pixel_data[159][9] = 0;
        pixel_data[159][10] = 0;
        pixel_data[159][11] = 0;
        pixel_data[159][12] = 0;
        pixel_data[159][13] = 0;
        pixel_data[159][14] = 0;
        pixel_data[159][15] = 0;
        pixel_data[159][16] = 0;
        pixel_data[159][17] = 13;
        pixel_data[159][18] = 11;
        pixel_data[159][19] = 11;
        pixel_data[159][20] = 8;
        pixel_data[159][21] = 5;
        pixel_data[159][22] = 1;
        pixel_data[159][23] = 1;
        pixel_data[159][24] = 1;
        pixel_data[159][25] = 1;
        pixel_data[159][26] = 1;
        pixel_data[159][27] = 1;
        pixel_data[159][28] = 1;
        pixel_data[159][29] = 1;
        pixel_data[159][30] = 1;
        pixel_data[159][31] = 1;
        pixel_data[159][32] = 1;
        pixel_data[159][33] = 1;
        pixel_data[159][34] = 1;
        pixel_data[159][35] = 1;
        pixel_data[159][36] = 1;
        pixel_data[159][37] = 1;
        pixel_data[159][38] = 1;
        pixel_data[159][39] = 1;
        pixel_data[159][40] = 1;
        pixel_data[159][41] = 1;
        pixel_data[159][42] = 1;
        pixel_data[159][43] = 1;
        pixel_data[159][44] = 1;
        pixel_data[159][45] = 1;
        pixel_data[159][46] = 1;
        pixel_data[159][47] = 1;
        pixel_data[159][48] = 1;
        pixel_data[159][49] = 1;
        pixel_data[159][50] = 1;
        pixel_data[159][51] = 1;
        pixel_data[159][52] = 1;
        pixel_data[159][53] = 1;
        pixel_data[159][54] = 1;
        pixel_data[159][55] = 1;
        pixel_data[159][56] = 1;
        pixel_data[159][57] = 1;
        pixel_data[159][58] = 1;
        pixel_data[159][59] = 1;
        pixel_data[159][60] = 1;
        pixel_data[159][61] = 1;
        pixel_data[159][62] = 1;
        pixel_data[159][63] = 1;
        pixel_data[159][64] = 1;
        pixel_data[159][65] = 1;
        pixel_data[159][66] = 1;
        pixel_data[159][67] = 1;
        pixel_data[159][68] = 1;
        pixel_data[159][69] = 1;
        pixel_data[159][70] = 1;
        pixel_data[159][71] = 1;
        pixel_data[159][72] = 1;
        pixel_data[159][73] = 1;
        pixel_data[159][74] = 1;
        pixel_data[159][75] = 1;
        pixel_data[159][76] = 1;
        pixel_data[159][77] = 1;
        pixel_data[159][78] = 1;
        pixel_data[159][79] = 1;
        pixel_data[159][80] = 1;
        pixel_data[159][81] = 1;
        pixel_data[159][82] = 1;
        pixel_data[159][83] = 1;
        pixel_data[159][84] = 1;
        pixel_data[159][85] = 1;
        pixel_data[159][86] = 1;
        pixel_data[159][87] = 1;
        pixel_data[159][88] = 1;
        pixel_data[159][89] = 1;
        pixel_data[159][90] = 1;
        pixel_data[159][91] = 1;
        pixel_data[159][92] = 1;
        pixel_data[159][93] = 1;
        pixel_data[159][94] = 1;
        pixel_data[159][95] = 1;
        pixel_data[159][96] = 6;
        pixel_data[159][97] = 8;
        pixel_data[159][98] = 10;
        pixel_data[159][99] = 12;
        pixel_data[159][100] = 13;
        pixel_data[159][101] = 13;
        pixel_data[159][102] = 13;
        pixel_data[159][103] = 13;
        pixel_data[159][104] = 13;
        pixel_data[159][105] = 13;
        pixel_data[159][106] = 13;
        pixel_data[159][107] = 13;
        pixel_data[159][108] = 12;
        pixel_data[159][109] = 12;
        pixel_data[159][110] = 9;
        pixel_data[159][111] = 6;
        pixel_data[159][112] = 1;
        pixel_data[159][113] = 1;
        pixel_data[159][114] = 1;
        pixel_data[159][115] = 1;
        pixel_data[159][116] = 1;
        pixel_data[159][117] = 1;
        pixel_data[159][118] = 1;
        pixel_data[159][119] = 1;
        pixel_data[159][120] = 1;
        pixel_data[159][121] = 1;
        pixel_data[159][122] = 1;
        pixel_data[159][123] = 1;
        pixel_data[159][124] = 1;
        pixel_data[159][125] = 1;
        pixel_data[159][126] = 1;
        pixel_data[159][127] = 1;
        pixel_data[159][128] = 1;
        pixel_data[159][129] = 1;
        pixel_data[159][130] = 1;
        pixel_data[159][131] = 1;
        pixel_data[159][132] = 1;
        pixel_data[159][133] = 1;
        pixel_data[159][134] = 4;
        pixel_data[159][135] = 6;
        pixel_data[159][136] = 7;
        pixel_data[159][137] = 8;
        pixel_data[159][138] = 9;
        pixel_data[159][139] = 8;
        pixel_data[159][140] = 7;
        pixel_data[159][141] = 6;
        pixel_data[159][142] = 4;
        pixel_data[159][143] = 1;
        pixel_data[159][144] = 1;
        pixel_data[159][145] = 1;
        pixel_data[159][146] = 1;
        pixel_data[159][147] = 1;
        pixel_data[159][148] = 1;
        pixel_data[159][149] = 1;
        pixel_data[159][150] = 1;
        pixel_data[159][151] = 1;
        pixel_data[159][152] = 1;
        pixel_data[159][153] = 1;
        pixel_data[159][154] = 1;
        pixel_data[159][155] = 1;
        pixel_data[159][156] = 1;
        pixel_data[159][157] = 1;
        pixel_data[159][158] = 1;
        pixel_data[159][159] = 1;
        pixel_data[159][160] = 1;
        pixel_data[159][161] = 1;
        pixel_data[159][162] = 1;
        pixel_data[159][163] = 1;
        pixel_data[159][164] = 1;
        pixel_data[159][165] = 1;
        pixel_data[159][166] = 1;
        pixel_data[159][167] = 1;
        pixel_data[159][168] = 1;
        pixel_data[159][169] = 1;
        pixel_data[159][170] = 7;
        pixel_data[159][171] = 9;
        pixel_data[159][172] = 11;
        pixel_data[159][173] = 11;
        pixel_data[159][174] = 0;
        pixel_data[159][175] = 0;
        pixel_data[159][176] = 0;
        pixel_data[159][177] = 0;
        pixel_data[159][178] = 0;
        pixel_data[159][179] = 0;
        pixel_data[159][180] = 0;
        pixel_data[159][181] = 0;
        pixel_data[159][182] = 0;
        pixel_data[159][183] = 0;
        pixel_data[159][184] = 0;
        pixel_data[159][185] = 0;
        pixel_data[159][186] = 0;
        pixel_data[159][187] = 0;
        pixel_data[159][188] = 0;
        pixel_data[159][189] = 0;
        pixel_data[159][190] = 0;
        pixel_data[159][191] = 0;
        pixel_data[159][192] = 0;
        pixel_data[159][193] = 0;
        pixel_data[159][194] = 0;
        pixel_data[159][195] = 0;
        pixel_data[159][196] = 0;
        pixel_data[159][197] = 0;
        pixel_data[159][198] = 0;
        pixel_data[159][199] = 0; // y=159
        pixel_data[160][0] = 0;
        pixel_data[160][1] = 0;
        pixel_data[160][2] = 0;
        pixel_data[160][3] = 0;
        pixel_data[160][4] = 0;
        pixel_data[160][5] = 0;
        pixel_data[160][6] = 0;
        pixel_data[160][7] = 0;
        pixel_data[160][8] = 0;
        pixel_data[160][9] = 0;
        pixel_data[160][10] = 0;
        pixel_data[160][11] = 0;
        pixel_data[160][12] = 0;
        pixel_data[160][13] = 0;
        pixel_data[160][14] = 0;
        pixel_data[160][15] = 0;
        pixel_data[160][16] = 0;
        pixel_data[160][17] = 11;
        pixel_data[160][18] = 11;
        pixel_data[160][19] = 8;
        pixel_data[160][20] = 5;
        pixel_data[160][21] = 1;
        pixel_data[160][22] = 1;
        pixel_data[160][23] = 1;
        pixel_data[160][24] = 1;
        pixel_data[160][25] = 1;
        pixel_data[160][26] = 1;
        pixel_data[160][27] = 1;
        pixel_data[160][28] = 1;
        pixel_data[160][29] = 1;
        pixel_data[160][30] = 1;
        pixel_data[160][31] = 1;
        pixel_data[160][32] = 1;
        pixel_data[160][33] = 1;
        pixel_data[160][34] = 1;
        pixel_data[160][35] = 1;
        pixel_data[160][36] = 1;
        pixel_data[160][37] = 1;
        pixel_data[160][38] = 1;
        pixel_data[160][39] = 1;
        pixel_data[160][40] = 1;
        pixel_data[160][41] = 1;
        pixel_data[160][42] = 1;
        pixel_data[160][43] = 1;
        pixel_data[160][44] = 1;
        pixel_data[160][45] = 1;
        pixel_data[160][46] = 1;
        pixel_data[160][47] = 1;
        pixel_data[160][48] = 1;
        pixel_data[160][49] = 1;
        pixel_data[160][50] = 1;
        pixel_data[160][51] = 1;
        pixel_data[160][52] = 1;
        pixel_data[160][53] = 1;
        pixel_data[160][54] = 1;
        pixel_data[160][55] = 1;
        pixel_data[160][56] = 1;
        pixel_data[160][57] = 1;
        pixel_data[160][58] = 1;
        pixel_data[160][59] = 1;
        pixel_data[160][60] = 1;
        pixel_data[160][61] = 1;
        pixel_data[160][62] = 1;
        pixel_data[160][63] = 1;
        pixel_data[160][64] = 1;
        pixel_data[160][65] = 1;
        pixel_data[160][66] = 1;
        pixel_data[160][67] = 1;
        pixel_data[160][68] = 1;
        pixel_data[160][69] = 1;
        pixel_data[160][70] = 1;
        pixel_data[160][71] = 1;
        pixel_data[160][72] = 1;
        pixel_data[160][73] = 1;
        pixel_data[160][74] = 1;
        pixel_data[160][75] = 1;
        pixel_data[160][76] = 1;
        pixel_data[160][77] = 1;
        pixel_data[160][78] = 1;
        pixel_data[160][79] = 1;
        pixel_data[160][80] = 1;
        pixel_data[160][81] = 1;
        pixel_data[160][82] = 1;
        pixel_data[160][83] = 1;
        pixel_data[160][84] = 1;
        pixel_data[160][85] = 1;
        pixel_data[160][86] = 1;
        pixel_data[160][87] = 1;
        pixel_data[160][88] = 1;
        pixel_data[160][89] = 1;
        pixel_data[160][90] = 1;
        pixel_data[160][91] = 1;
        pixel_data[160][92] = 4;
        pixel_data[160][93] = 7;
        pixel_data[160][94] = 10;
        pixel_data[160][95] = 12;
        pixel_data[160][96] = 13;
        pixel_data[160][97] = 13;
        pixel_data[160][98] = 13;
        pixel_data[160][99] = 13;
        pixel_data[160][100] = 13;
        pixel_data[160][101] = 13;
        pixel_data[160][102] = 13;
        pixel_data[160][103] = 13;
        pixel_data[160][104] = 13;
        pixel_data[160][105] = 13;
        pixel_data[160][106] = 13;
        pixel_data[160][107] = 13;
        pixel_data[160][108] = 13;
        pixel_data[160][109] = 13;
        pixel_data[160][110] = 13;
        pixel_data[160][111] = 13;
        pixel_data[160][112] = 12;
        pixel_data[160][113] = 8;
        pixel_data[160][114] = 4;
        pixel_data[160][115] = 1;
        pixel_data[160][116] = 1;
        pixel_data[160][117] = 1;
        pixel_data[160][118] = 1;
        pixel_data[160][119] = 1;
        pixel_data[160][120] = 1;
        pixel_data[160][121] = 1;
        pixel_data[160][122] = 1;
        pixel_data[160][123] = 1;
        pixel_data[160][124] = 1;
        pixel_data[160][125] = 1;
        pixel_data[160][126] = 1;
        pixel_data[160][127] = 1;
        pixel_data[160][128] = 1;
        pixel_data[160][129] = 1;
        pixel_data[160][130] = 1;
        pixel_data[160][131] = 5;
        pixel_data[160][132] = 9;
        pixel_data[160][133] = 12;
        pixel_data[160][134] = 13;
        pixel_data[160][135] = 13;
        pixel_data[160][136] = 13;
        pixel_data[160][137] = 13;
        pixel_data[160][138] = 13;
        pixel_data[160][139] = 13;
        pixel_data[160][140] = 13;
        pixel_data[160][141] = 13;
        pixel_data[160][142] = 13;
        pixel_data[160][143] = 13;
        pixel_data[160][144] = 13;
        pixel_data[160][145] = 13;
        pixel_data[160][146] = 9;
        pixel_data[160][147] = 5;
        pixel_data[160][148] = 1;
        pixel_data[160][149] = 1;
        pixel_data[160][150] = 1;
        pixel_data[160][151] = 1;
        pixel_data[160][152] = 1;
        pixel_data[160][153] = 1;
        pixel_data[160][154] = 1;
        pixel_data[160][155] = 1;
        pixel_data[160][156] = 1;
        pixel_data[160][157] = 1;
        pixel_data[160][158] = 1;
        pixel_data[160][159] = 1;
        pixel_data[160][160] = 1;
        pixel_data[160][161] = 1;
        pixel_data[160][162] = 1;
        pixel_data[160][163] = 1;
        pixel_data[160][164] = 1;
        pixel_data[160][165] = 1;
        pixel_data[160][166] = 1;
        pixel_data[160][167] = 1;
        pixel_data[160][168] = 1;
        pixel_data[160][169] = 1;
        pixel_data[160][170] = 1;
        pixel_data[160][171] = 5;
        pixel_data[160][172] = 8;
        pixel_data[160][173] = 11;
        pixel_data[160][174] = 11;
        pixel_data[160][175] = 0;
        pixel_data[160][176] = 0;
        pixel_data[160][177] = 0;
        pixel_data[160][178] = 0;
        pixel_data[160][179] = 0;
        pixel_data[160][180] = 0;
        pixel_data[160][181] = 0;
        pixel_data[160][182] = 0;
        pixel_data[160][183] = 0;
        pixel_data[160][184] = 0;
        pixel_data[160][185] = 0;
        pixel_data[160][186] = 0;
        pixel_data[160][187] = 0;
        pixel_data[160][188] = 0;
        pixel_data[160][189] = 0;
        pixel_data[160][190] = 0;
        pixel_data[160][191] = 0;
        pixel_data[160][192] = 0;
        pixel_data[160][193] = 0;
        pixel_data[160][194] = 0;
        pixel_data[160][195] = 0;
        pixel_data[160][196] = 0;
        pixel_data[160][197] = 0;
        pixel_data[160][198] = 0;
        pixel_data[160][199] = 0; // y=160
        pixel_data[161][0] = 0;
        pixel_data[161][1] = 0;
        pixel_data[161][2] = 0;
        pixel_data[161][3] = 0;
        pixel_data[161][4] = 0;
        pixel_data[161][5] = 0;
        pixel_data[161][6] = 0;
        pixel_data[161][7] = 0;
        pixel_data[161][8] = 0;
        pixel_data[161][9] = 0;
        pixel_data[161][10] = 0;
        pixel_data[161][11] = 0;
        pixel_data[161][12] = 0;
        pixel_data[161][13] = 0;
        pixel_data[161][14] = 0;
        pixel_data[161][15] = 0;
        pixel_data[161][16] = 11;
        pixel_data[161][17] = 11;
        pixel_data[161][18] = 8;
        pixel_data[161][19] = 5;
        pixel_data[161][20] = 1;
        pixel_data[161][21] = 1;
        pixel_data[161][22] = 1;
        pixel_data[161][23] = 1;
        pixel_data[161][24] = 1;
        pixel_data[161][25] = 1;
        pixel_data[161][26] = 1;
        pixel_data[161][27] = 1;
        pixel_data[161][28] = 1;
        pixel_data[161][29] = 1;
        pixel_data[161][30] = 1;
        pixel_data[161][31] = 1;
        pixel_data[161][32] = 1;
        pixel_data[161][33] = 1;
        pixel_data[161][34] = 1;
        pixel_data[161][35] = 1;
        pixel_data[161][36] = 1;
        pixel_data[161][37] = 1;
        pixel_data[161][38] = 1;
        pixel_data[161][39] = 1;
        pixel_data[161][40] = 1;
        pixel_data[161][41] = 1;
        pixel_data[161][42] = 1;
        pixel_data[161][43] = 1;
        pixel_data[161][44] = 1;
        pixel_data[161][45] = 1;
        pixel_data[161][46] = 1;
        pixel_data[161][47] = 1;
        pixel_data[161][48] = 1;
        pixel_data[161][49] = 1;
        pixel_data[161][50] = 1;
        pixel_data[161][51] = 1;
        pixel_data[161][52] = 1;
        pixel_data[161][53] = 1;
        pixel_data[161][54] = 1;
        pixel_data[161][55] = 1;
        pixel_data[161][56] = 1;
        pixel_data[161][57] = 1;
        pixel_data[161][58] = 1;
        pixel_data[161][59] = 1;
        pixel_data[161][60] = 1;
        pixel_data[161][61] = 1;
        pixel_data[161][62] = 1;
        pixel_data[161][63] = 1;
        pixel_data[161][64] = 1;
        pixel_data[161][65] = 1;
        pixel_data[161][66] = 1;
        pixel_data[161][67] = 1;
        pixel_data[161][68] = 1;
        pixel_data[161][69] = 1;
        pixel_data[161][70] = 1;
        pixel_data[161][71] = 1;
        pixel_data[161][72] = 1;
        pixel_data[161][73] = 1;
        pixel_data[161][74] = 1;
        pixel_data[161][75] = 1;
        pixel_data[161][76] = 1;
        pixel_data[161][77] = 1;
        pixel_data[161][78] = 1;
        pixel_data[161][79] = 1;
        pixel_data[161][80] = 1;
        pixel_data[161][81] = 1;
        pixel_data[161][82] = 1;
        pixel_data[161][83] = 1;
        pixel_data[161][84] = 1;
        pixel_data[161][85] = 1;
        pixel_data[161][86] = 1;
        pixel_data[161][87] = 1;
        pixel_data[161][88] = 1;
        pixel_data[161][89] = 1;
        pixel_data[161][90] = 6;
        pixel_data[161][91] = 9;
        pixel_data[161][92] = 12;
        pixel_data[161][93] = 13;
        pixel_data[161][94] = 13;
        pixel_data[161][95] = 13;
        pixel_data[161][96] = 13;
        pixel_data[161][97] = 13;
        pixel_data[161][98] = 13;
        pixel_data[161][99] = 13;
        pixel_data[161][100] = 13;
        pixel_data[161][101] = 13;
        pixel_data[161][102] = 13;
        pixel_data[161][103] = 13;
        pixel_data[161][104] = 13;
        pixel_data[161][105] = 13;
        pixel_data[161][106] = 13;
        pixel_data[161][107] = 13;
        pixel_data[161][108] = 13;
        pixel_data[161][109] = 13;
        pixel_data[161][110] = 13;
        pixel_data[161][111] = 13;
        pixel_data[161][112] = 13;
        pixel_data[161][113] = 13;
        pixel_data[161][114] = 10;
        pixel_data[161][115] = 6;
        pixel_data[161][116] = 1;
        pixel_data[161][117] = 1;
        pixel_data[161][118] = 1;
        pixel_data[161][119] = 1;
        pixel_data[161][120] = 1;
        pixel_data[161][121] = 1;
        pixel_data[161][122] = 1;
        pixel_data[161][123] = 1;
        pixel_data[161][124] = 1;
        pixel_data[161][125] = 1;
        pixel_data[161][126] = 1;
        pixel_data[161][127] = 1;
        pixel_data[161][128] = 1;
        pixel_data[161][129] = 5;
        pixel_data[161][130] = 9;
        pixel_data[161][131] = 12;
        pixel_data[161][132] = 13;
        pixel_data[161][133] = 13;
        pixel_data[161][134] = 13;
        pixel_data[161][135] = 13;
        pixel_data[161][136] = 13;
        pixel_data[161][137] = 13;
        pixel_data[161][138] = 13;
        pixel_data[161][139] = 13;
        pixel_data[161][140] = 13;
        pixel_data[161][141] = 13;
        pixel_data[161][142] = 13;
        pixel_data[161][143] = 13;
        pixel_data[161][144] = 13;
        pixel_data[161][145] = 13;
        pixel_data[161][146] = 13;
        pixel_data[161][147] = 13;
        pixel_data[161][148] = 12;
        pixel_data[161][149] = 7;
        pixel_data[161][150] = 2;
        pixel_data[161][151] = 1;
        pixel_data[161][152] = 1;
        pixel_data[161][153] = 1;
        pixel_data[161][154] = 1;
        pixel_data[161][155] = 1;
        pixel_data[161][156] = 1;
        pixel_data[161][157] = 1;
        pixel_data[161][158] = 1;
        pixel_data[161][159] = 1;
        pixel_data[161][160] = 1;
        pixel_data[161][161] = 1;
        pixel_data[161][162] = 1;
        pixel_data[161][163] = 1;
        pixel_data[161][164] = 1;
        pixel_data[161][165] = 1;
        pixel_data[161][166] = 1;
        pixel_data[161][167] = 1;
        pixel_data[161][168] = 1;
        pixel_data[161][169] = 1;
        pixel_data[161][170] = 1;
        pixel_data[161][171] = 1;
        pixel_data[161][172] = 4;
        pixel_data[161][173] = 7;
        pixel_data[161][174] = 9;
        pixel_data[161][175] = 11;
        pixel_data[161][176] = 13;
        pixel_data[161][177] = 0;
        pixel_data[161][178] = 0;
        pixel_data[161][179] = 0;
        pixel_data[161][180] = 0;
        pixel_data[161][181] = 0;
        pixel_data[161][182] = 0;
        pixel_data[161][183] = 0;
        pixel_data[161][184] = 0;
        pixel_data[161][185] = 0;
        pixel_data[161][186] = 0;
        pixel_data[161][187] = 0;
        pixel_data[161][188] = 0;
        pixel_data[161][189] = 0;
        pixel_data[161][190] = 0;
        pixel_data[161][191] = 0;
        pixel_data[161][192] = 0;
        pixel_data[161][193] = 0;
        pixel_data[161][194] = 0;
        pixel_data[161][195] = 0;
        pixel_data[161][196] = 0;
        pixel_data[161][197] = 0;
        pixel_data[161][198] = 0;
        pixel_data[161][199] = 0; // y=161
        pixel_data[162][0] = 0;
        pixel_data[162][1] = 0;
        pixel_data[162][2] = 0;
        pixel_data[162][3] = 0;
        pixel_data[162][4] = 0;
        pixel_data[162][5] = 0;
        pixel_data[162][6] = 0;
        pixel_data[162][7] = 0;
        pixel_data[162][8] = 0;
        pixel_data[162][9] = 0;
        pixel_data[162][10] = 0;
        pixel_data[162][11] = 0;
        pixel_data[162][12] = 0;
        pixel_data[162][13] = 0;
        pixel_data[162][14] = 10;
        pixel_data[162][15] = 11;
        pixel_data[162][16] = 9;
        pixel_data[162][17] = 7;
        pixel_data[162][18] = 1;
        pixel_data[162][19] = 1;
        pixel_data[162][20] = 1;
        pixel_data[162][21] = 1;
        pixel_data[162][22] = 1;
        pixel_data[162][23] = 1;
        pixel_data[162][24] = 1;
        pixel_data[162][25] = 1;
        pixel_data[162][26] = 1;
        pixel_data[162][27] = 1;
        pixel_data[162][28] = 1;
        pixel_data[162][29] = 1;
        pixel_data[162][30] = 1;
        pixel_data[162][31] = 1;
        pixel_data[162][32] = 1;
        pixel_data[162][33] = 1;
        pixel_data[162][34] = 1;
        pixel_data[162][35] = 1;
        pixel_data[162][36] = 1;
        pixel_data[162][37] = 1;
        pixel_data[162][38] = 1;
        pixel_data[162][39] = 1;
        pixel_data[162][40] = 1;
        pixel_data[162][41] = 1;
        pixel_data[162][42] = 1;
        pixel_data[162][43] = 1;
        pixel_data[162][44] = 1;
        pixel_data[162][45] = 1;
        pixel_data[162][46] = 1;
        pixel_data[162][47] = 1;
        pixel_data[162][48] = 1;
        pixel_data[162][49] = 1;
        pixel_data[162][50] = 1;
        pixel_data[162][51] = 1;
        pixel_data[162][52] = 1;
        pixel_data[162][53] = 1;
        pixel_data[162][54] = 1;
        pixel_data[162][55] = 1;
        pixel_data[162][56] = 1;
        pixel_data[162][57] = 1;
        pixel_data[162][58] = 1;
        pixel_data[162][59] = 1;
        pixel_data[162][60] = 1;
        pixel_data[162][61] = 1;
        pixel_data[162][62] = 1;
        pixel_data[162][63] = 1;
        pixel_data[162][64] = 1;
        pixel_data[162][65] = 1;
        pixel_data[162][66] = 1;
        pixel_data[162][67] = 1;
        pixel_data[162][68] = 1;
        pixel_data[162][69] = 1;
        pixel_data[162][70] = 1;
        pixel_data[162][71] = 1;
        pixel_data[162][72] = 1;
        pixel_data[162][73] = 1;
        pixel_data[162][74] = 1;
        pixel_data[162][75] = 1;
        pixel_data[162][76] = 1;
        pixel_data[162][77] = 1;
        pixel_data[162][78] = 1;
        pixel_data[162][79] = 1;
        pixel_data[162][80] = 1;
        pixel_data[162][81] = 1;
        pixel_data[162][82] = 1;
        pixel_data[162][83] = 1;
        pixel_data[162][84] = 1;
        pixel_data[162][85] = 1;
        pixel_data[162][86] = 1;
        pixel_data[162][87] = 4;
        pixel_data[162][88] = 8;
        pixel_data[162][89] = 12;
        pixel_data[162][90] = 13;
        pixel_data[162][91] = 13;
        pixel_data[162][92] = 13;
        pixel_data[162][93] = 13;
        pixel_data[162][94] = 13;
        pixel_data[162][95] = 13;
        pixel_data[162][96] = 13;
        pixel_data[162][97] = 13;
        pixel_data[162][98] = 13;
        pixel_data[162][99] = 13;
        pixel_data[162][100] = 13;
        pixel_data[162][101] = 13;
        pixel_data[162][102] = 13;
        pixel_data[162][103] = 13;
        pixel_data[162][104] = 13;
        pixel_data[162][105] = 13;
        pixel_data[162][106] = 13;
        pixel_data[162][107] = 13;
        pixel_data[162][108] = 13;
        pixel_data[162][109] = 13;
        pixel_data[162][110] = 13;
        pixel_data[162][111] = 13;
        pixel_data[162][112] = 13;
        pixel_data[162][113] = 13;
        pixel_data[162][114] = 13;
        pixel_data[162][115] = 10;
        pixel_data[162][116] = 5;
        pixel_data[162][117] = 1;
        pixel_data[162][118] = 1;
        pixel_data[162][119] = 1;
        pixel_data[162][120] = 1;
        pixel_data[162][121] = 1;
        pixel_data[162][122] = 1;
        pixel_data[162][123] = 1;
        pixel_data[162][124] = 1;
        pixel_data[162][125] = 1;
        pixel_data[162][126] = 1;
        pixel_data[162][127] = 1;
        pixel_data[162][128] = 6;
        pixel_data[162][129] = 10;
        pixel_data[162][130] = 13;
        pixel_data[162][131] = 13;
        pixel_data[162][132] = 13;
        pixel_data[162][133] = 13;
        pixel_data[162][134] = 13;
        pixel_data[162][135] = 13;
        pixel_data[162][136] = 13;
        pixel_data[162][137] = 13;
        pixel_data[162][138] = 13;
        pixel_data[162][139] = 13;
        pixel_data[162][140] = 13;
        pixel_data[162][141] = 13;
        pixel_data[162][142] = 13;
        pixel_data[162][143] = 13;
        pixel_data[162][144] = 13;
        pixel_data[162][145] = 13;
        pixel_data[162][146] = 13;
        pixel_data[162][147] = 13;
        pixel_data[162][148] = 13;
        pixel_data[162][149] = 13;
        pixel_data[162][150] = 13;
        pixel_data[162][151] = 10;
        pixel_data[162][152] = 4;
        pixel_data[162][153] = 1;
        pixel_data[162][154] = 1;
        pixel_data[162][155] = 1;
        pixel_data[162][156] = 1;
        pixel_data[162][157] = 1;
        pixel_data[162][158] = 1;
        pixel_data[162][159] = 1;
        pixel_data[162][160] = 1;
        pixel_data[162][161] = 1;
        pixel_data[162][162] = 1;
        pixel_data[162][163] = 1;
        pixel_data[162][164] = 1;
        pixel_data[162][165] = 1;
        pixel_data[162][166] = 1;
        pixel_data[162][167] = 1;
        pixel_data[162][168] = 1;
        pixel_data[162][169] = 1;
        pixel_data[162][170] = 1;
        pixel_data[162][171] = 1;
        pixel_data[162][172] = 1;
        pixel_data[162][173] = 1;
        pixel_data[162][174] = 6;
        pixel_data[162][175] = 9;
        pixel_data[162][176] = 11;
        pixel_data[162][177] = 11;
        pixel_data[162][178] = 0;
        pixel_data[162][179] = 0;
        pixel_data[162][180] = 0;
        pixel_data[162][181] = 0;
        pixel_data[162][182] = 0;
        pixel_data[162][183] = 0;
        pixel_data[162][184] = 0;
        pixel_data[162][185] = 0;
        pixel_data[162][186] = 0;
        pixel_data[162][187] = 0;
        pixel_data[162][188] = 0;
        pixel_data[162][189] = 0;
        pixel_data[162][190] = 0;
        pixel_data[162][191] = 0;
        pixel_data[162][192] = 0;
        pixel_data[162][193] = 0;
        pixel_data[162][194] = 0;
        pixel_data[162][195] = 0;
        pixel_data[162][196] = 0;
        pixel_data[162][197] = 0;
        pixel_data[162][198] = 0;
        pixel_data[162][199] = 0; // y=162
        pixel_data[163][0] = 0;
        pixel_data[163][1] = 0;
        pixel_data[163][2] = 0;
        pixel_data[163][3] = 0;
        pixel_data[163][4] = 0;
        pixel_data[163][5] = 0;
        pixel_data[163][6] = 0;
        pixel_data[163][7] = 0;
        pixel_data[163][8] = 0;
        pixel_data[163][9] = 0;
        pixel_data[163][10] = 0;
        pixel_data[163][11] = 0;
        pixel_data[163][12] = 0;
        pixel_data[163][13] = 10;
        pixel_data[163][14] = 11;
        pixel_data[163][15] = 9;
        pixel_data[163][16] = 7;
        pixel_data[163][17] = 4;
        pixel_data[163][18] = 1;
        pixel_data[163][19] = 1;
        pixel_data[163][20] = 1;
        pixel_data[163][21] = 1;
        pixel_data[163][22] = 1;
        pixel_data[163][23] = 1;
        pixel_data[163][24] = 1;
        pixel_data[163][25] = 1;
        pixel_data[163][26] = 1;
        pixel_data[163][27] = 1;
        pixel_data[163][28] = 1;
        pixel_data[163][29] = 1;
        pixel_data[163][30] = 1;
        pixel_data[163][31] = 1;
        pixel_data[163][32] = 1;
        pixel_data[163][33] = 1;
        pixel_data[163][34] = 1;
        pixel_data[163][35] = 1;
        pixel_data[163][36] = 1;
        pixel_data[163][37] = 1;
        pixel_data[163][38] = 1;
        pixel_data[163][39] = 1;
        pixel_data[163][40] = 1;
        pixel_data[163][41] = 1;
        pixel_data[163][42] = 1;
        pixel_data[163][43] = 1;
        pixel_data[163][44] = 1;
        pixel_data[163][45] = 1;
        pixel_data[163][46] = 1;
        pixel_data[163][47] = 1;
        pixel_data[163][48] = 1;
        pixel_data[163][49] = 1;
        pixel_data[163][50] = 1;
        pixel_data[163][51] = 1;
        pixel_data[163][52] = 1;
        pixel_data[163][53] = 1;
        pixel_data[163][54] = 1;
        pixel_data[163][55] = 1;
        pixel_data[163][56] = 1;
        pixel_data[163][57] = 1;
        pixel_data[163][58] = 1;
        pixel_data[163][59] = 1;
        pixel_data[163][60] = 1;
        pixel_data[163][61] = 1;
        pixel_data[163][62] = 1;
        pixel_data[163][63] = 1;
        pixel_data[163][64] = 1;
        pixel_data[163][65] = 1;
        pixel_data[163][66] = 1;
        pixel_data[163][67] = 1;
        pixel_data[163][68] = 1;
        pixel_data[163][69] = 1;
        pixel_data[163][70] = 1;
        pixel_data[163][71] = 1;
        pixel_data[163][72] = 1;
        pixel_data[163][73] = 1;
        pixel_data[163][74] = 1;
        pixel_data[163][75] = 1;
        pixel_data[163][76] = 1;
        pixel_data[163][77] = 1;
        pixel_data[163][78] = 1;
        pixel_data[163][79] = 1;
        pixel_data[163][80] = 1;
        pixel_data[163][81] = 1;
        pixel_data[163][82] = 1;
        pixel_data[163][83] = 1;
        pixel_data[163][84] = 1;
        pixel_data[163][85] = 1;
        pixel_data[163][86] = 5;
        pixel_data[163][87] = 10;
        pixel_data[163][88] = 13;
        pixel_data[163][89] = 13;
        pixel_data[163][90] = 13;
        pixel_data[163][91] = 13;
        pixel_data[163][92] = 13;
        pixel_data[163][93] = 13;
        pixel_data[163][94] = 13;
        pixel_data[163][95] = 13;
        pixel_data[163][96] = 13;
        pixel_data[163][97] = 13;
        pixel_data[163][98] = 13;
        pixel_data[163][99] = 13;
        pixel_data[163][100] = 13;
        pixel_data[163][101] = 13;
        pixel_data[163][102] = 13;
        pixel_data[163][103] = 13;
        pixel_data[163][104] = 13;
        pixel_data[163][105] = 13;
        pixel_data[163][106] = 13;
        pixel_data[163][107] = 13;
        pixel_data[163][108] = 13;
        pixel_data[163][109] = 13;
        pixel_data[163][110] = 13;
        pixel_data[163][111] = 13;
        pixel_data[163][112] = 13;
        pixel_data[163][113] = 13;
        pixel_data[163][114] = 13;
        pixel_data[163][115] = 12;
        pixel_data[163][116] = 7;
        pixel_data[163][117] = 1;
        pixel_data[163][118] = 1;
        pixel_data[163][119] = 1;
        pixel_data[163][120] = 1;
        pixel_data[163][121] = 1;
        pixel_data[163][122] = 1;
        pixel_data[163][123] = 1;
        pixel_data[163][124] = 1;
        pixel_data[163][125] = 1;
        pixel_data[163][126] = 1;
        pixel_data[163][127] = 1;
        pixel_data[163][128] = 5;
        pixel_data[163][129] = 12;
        pixel_data[163][130] = 13;
        pixel_data[163][131] = 13;
        pixel_data[163][132] = 13;
        pixel_data[163][133] = 13;
        pixel_data[163][134] = 13;
        pixel_data[163][135] = 13;
        pixel_data[163][136] = 13;
        pixel_data[163][137] = 13;
        pixel_data[163][138] = 13;
        pixel_data[163][139] = 13;
        pixel_data[163][140] = 13;
        pixel_data[163][141] = 13;
        pixel_data[163][142] = 13;
        pixel_data[163][143] = 13;
        pixel_data[163][144] = 13;
        pixel_data[163][145] = 13;
        pixel_data[163][146] = 13;
        pixel_data[163][147] = 13;
        pixel_data[163][148] = 13;
        pixel_data[163][149] = 13;
        pixel_data[163][150] = 13;
        pixel_data[163][151] = 13;
        pixel_data[163][152] = 10;
        pixel_data[163][153] = 4;
        pixel_data[163][154] = 1;
        pixel_data[163][155] = 1;
        pixel_data[163][156] = 1;
        pixel_data[163][157] = 1;
        pixel_data[163][158] = 1;
        pixel_data[163][159] = 1;
        pixel_data[163][160] = 1;
        pixel_data[163][161] = 1;
        pixel_data[163][162] = 1;
        pixel_data[163][163] = 1;
        pixel_data[163][164] = 1;
        pixel_data[163][165] = 1;
        pixel_data[163][166] = 1;
        pixel_data[163][167] = 1;
        pixel_data[163][168] = 1;
        pixel_data[163][169] = 1;
        pixel_data[163][170] = 1;
        pixel_data[163][171] = 1;
        pixel_data[163][172] = 1;
        pixel_data[163][173] = 1;
        pixel_data[163][174] = 1;
        pixel_data[163][175] = 6;
        pixel_data[163][176] = 9;
        pixel_data[163][177] = 11;
        pixel_data[163][178] = 11;
        pixel_data[163][179] = 0;
        pixel_data[163][180] = 0;
        pixel_data[163][181] = 0;
        pixel_data[163][182] = 0;
        pixel_data[163][183] = 0;
        pixel_data[163][184] = 0;
        pixel_data[163][185] = 0;
        pixel_data[163][186] = 0;
        pixel_data[163][187] = 0;
        pixel_data[163][188] = 0;
        pixel_data[163][189] = 0;
        pixel_data[163][190] = 0;
        pixel_data[163][191] = 0;
        pixel_data[163][192] = 0;
        pixel_data[163][193] = 0;
        pixel_data[163][194] = 0;
        pixel_data[163][195] = 0;
        pixel_data[163][196] = 0;
        pixel_data[163][197] = 0;
        pixel_data[163][198] = 0;
        pixel_data[163][199] = 0; // y=163
        pixel_data[164][0] = 0;
        pixel_data[164][1] = 0;
        pixel_data[164][2] = 0;
        pixel_data[164][3] = 0;
        pixel_data[164][4] = 0;
        pixel_data[164][5] = 0;
        pixel_data[164][6] = 0;
        pixel_data[164][7] = 0;
        pixel_data[164][8] = 0;
        pixel_data[164][9] = 0;
        pixel_data[164][10] = 0;
        pixel_data[164][11] = 0;
        pixel_data[164][12] = 11;
        pixel_data[164][13] = 11;
        pixel_data[164][14] = 9;
        pixel_data[164][15] = 7;
        pixel_data[164][16] = 4;
        pixel_data[164][17] = 2;
        pixel_data[164][18] = 1;
        pixel_data[164][19] = 1;
        pixel_data[164][20] = 1;
        pixel_data[164][21] = 1;
        pixel_data[164][22] = 1;
        pixel_data[164][23] = 1;
        pixel_data[164][24] = 1;
        pixel_data[164][25] = 1;
        pixel_data[164][26] = 1;
        pixel_data[164][27] = 1;
        pixel_data[164][28] = 1;
        pixel_data[164][29] = 1;
        pixel_data[164][30] = 1;
        pixel_data[164][31] = 1;
        pixel_data[164][32] = 1;
        pixel_data[164][33] = 1;
        pixel_data[164][34] = 1;
        pixel_data[164][35] = 1;
        pixel_data[164][36] = 1;
        pixel_data[164][37] = 1;
        pixel_data[164][38] = 1;
        pixel_data[164][39] = 1;
        pixel_data[164][40] = 1;
        pixel_data[164][41] = 1;
        pixel_data[164][42] = 1;
        pixel_data[164][43] = 1;
        pixel_data[164][44] = 1;
        pixel_data[164][45] = 1;
        pixel_data[164][46] = 1;
        pixel_data[164][47] = 1;
        pixel_data[164][48] = 1;
        pixel_data[164][49] = 1;
        pixel_data[164][50] = 1;
        pixel_data[164][51] = 1;
        pixel_data[164][52] = 1;
        pixel_data[164][53] = 1;
        pixel_data[164][54] = 1;
        pixel_data[164][55] = 1;
        pixel_data[164][56] = 1;
        pixel_data[164][57] = 1;
        pixel_data[164][58] = 1;
        pixel_data[164][59] = 1;
        pixel_data[164][60] = 1;
        pixel_data[164][61] = 1;
        pixel_data[164][62] = 1;
        pixel_data[164][63] = 1;
        pixel_data[164][64] = 1;
        pixel_data[164][65] = 1;
        pixel_data[164][66] = 1;
        pixel_data[164][67] = 1;
        pixel_data[164][68] = 1;
        pixel_data[164][69] = 1;
        pixel_data[164][70] = 1;
        pixel_data[164][71] = 1;
        pixel_data[164][72] = 1;
        pixel_data[164][73] = 1;
        pixel_data[164][74] = 1;
        pixel_data[164][75] = 1;
        pixel_data[164][76] = 1;
        pixel_data[164][77] = 1;
        pixel_data[164][78] = 1;
        pixel_data[164][79] = 1;
        pixel_data[164][80] = 1;
        pixel_data[164][81] = 1;
        pixel_data[164][82] = 1;
        pixel_data[164][83] = 1;
        pixel_data[164][84] = 1;
        pixel_data[164][85] = 1;
        pixel_data[164][86] = 7;
        pixel_data[164][87] = 12;
        pixel_data[164][88] = 13;
        pixel_data[164][89] = 13;
        pixel_data[164][90] = 13;
        pixel_data[164][91] = 13;
        pixel_data[164][92] = 13;
        pixel_data[164][93] = 13;
        pixel_data[164][94] = 13;
        pixel_data[164][95] = 13;
        pixel_data[164][96] = 13;
        pixel_data[164][97] = 13;
        pixel_data[164][98] = 13;
        pixel_data[164][99] = 13;
        pixel_data[164][100] = 13;
        pixel_data[164][101] = 13;
        pixel_data[164][102] = 13;
        pixel_data[164][103] = 13;
        pixel_data[164][104] = 13;
        pixel_data[164][105] = 13;
        pixel_data[164][106] = 13;
        pixel_data[164][107] = 13;
        pixel_data[164][108] = 13;
        pixel_data[164][109] = 13;
        pixel_data[164][110] = 13;
        pixel_data[164][111] = 13;
        pixel_data[164][112] = 13;
        pixel_data[164][113] = 13;
        pixel_data[164][114] = 13;
        pixel_data[164][115] = 13;
        pixel_data[164][116] = 9;
        pixel_data[164][117] = 1;
        pixel_data[164][118] = 1;
        pixel_data[164][119] = 1;
        pixel_data[164][120] = 1;
        pixel_data[164][121] = 1;
        pixel_data[164][122] = 1;
        pixel_data[164][123] = 1;
        pixel_data[164][124] = 1;
        pixel_data[164][125] = 1;
        pixel_data[164][126] = 1;
        pixel_data[164][127] = 1;
        pixel_data[164][128] = 1;
        pixel_data[164][129] = 8;
        pixel_data[164][130] = 12;
        pixel_data[164][131] = 13;
        pixel_data[164][132] = 13;
        pixel_data[164][133] = 13;
        pixel_data[164][134] = 13;
        pixel_data[164][135] = 13;
        pixel_data[164][136] = 13;
        pixel_data[164][137] = 13;
        pixel_data[164][138] = 13;
        pixel_data[164][139] = 13;
        pixel_data[164][140] = 13;
        pixel_data[164][141] = 13;
        pixel_data[164][142] = 13;
        pixel_data[164][143] = 13;
        pixel_data[164][144] = 13;
        pixel_data[164][145] = 13;
        pixel_data[164][146] = 13;
        pixel_data[164][147] = 13;
        pixel_data[164][148] = 13;
        pixel_data[164][149] = 13;
        pixel_data[164][150] = 13;
        pixel_data[164][151] = 13;
        pixel_data[164][152] = 13;
        pixel_data[164][153] = 8;
        pixel_data[164][154] = 1;
        pixel_data[164][155] = 1;
        pixel_data[164][156] = 1;
        pixel_data[164][157] = 1;
        pixel_data[164][158] = 1;
        pixel_data[164][159] = 1;
        pixel_data[164][160] = 1;
        pixel_data[164][161] = 1;
        pixel_data[164][162] = 1;
        pixel_data[164][163] = 1;
        pixel_data[164][164] = 1;
        pixel_data[164][165] = 1;
        pixel_data[164][166] = 1;
        pixel_data[164][167] = 1;
        pixel_data[164][168] = 1;
        pixel_data[164][169] = 1;
        pixel_data[164][170] = 1;
        pixel_data[164][171] = 1;
        pixel_data[164][172] = 1;
        pixel_data[164][173] = 1;
        pixel_data[164][174] = 1;
        pixel_data[164][175] = 1;
        pixel_data[164][176] = 7;
        pixel_data[164][177] = 9;
        pixel_data[164][178] = 11;
        pixel_data[164][179] = 10;
        pixel_data[164][180] = 0;
        pixel_data[164][181] = 0;
        pixel_data[164][182] = 0;
        pixel_data[164][183] = 0;
        pixel_data[164][184] = 0;
        pixel_data[164][185] = 0;
        pixel_data[164][186] = 0;
        pixel_data[164][187] = 0;
        pixel_data[164][188] = 0;
        pixel_data[164][189] = 0;
        pixel_data[164][190] = 0;
        pixel_data[164][191] = 0;
        pixel_data[164][192] = 0;
        pixel_data[164][193] = 0;
        pixel_data[164][194] = 0;
        pixel_data[164][195] = 0;
        pixel_data[164][196] = 0;
        pixel_data[164][197] = 0;
        pixel_data[164][198] = 0;
        pixel_data[164][199] = 0; // y=164
        pixel_data[165][0] = 0;
        pixel_data[165][1] = 0;
        pixel_data[165][2] = 0;
        pixel_data[165][3] = 0;
        pixel_data[165][4] = 0;
        pixel_data[165][5] = 0;
        pixel_data[165][6] = 0;
        pixel_data[165][7] = 0;
        pixel_data[165][8] = 0;
        pixel_data[165][9] = 0;
        pixel_data[165][10] = 0;
        pixel_data[165][11] = 11;
        pixel_data[165][12] = 11;
        pixel_data[165][13] = 9;
        pixel_data[165][14] = 7;
        pixel_data[165][15] = 4;
        pixel_data[165][16] = 4;
        pixel_data[165][17] = 1;
        pixel_data[165][18] = 1;
        pixel_data[165][19] = 1;
        pixel_data[165][20] = 1;
        pixel_data[165][21] = 1;
        pixel_data[165][22] = 1;
        pixel_data[165][23] = 1;
        pixel_data[165][24] = 1;
        pixel_data[165][25] = 1;
        pixel_data[165][26] = 1;
        pixel_data[165][27] = 1;
        pixel_data[165][28] = 1;
        pixel_data[165][29] = 1;
        pixel_data[165][30] = 1;
        pixel_data[165][31] = 1;
        pixel_data[165][32] = 1;
        pixel_data[165][33] = 1;
        pixel_data[165][34] = 1;
        pixel_data[165][35] = 1;
        pixel_data[165][36] = 1;
        pixel_data[165][37] = 1;
        pixel_data[165][38] = 1;
        pixel_data[165][39] = 1;
        pixel_data[165][40] = 1;
        pixel_data[165][41] = 1;
        pixel_data[165][42] = 1;
        pixel_data[165][43] = 1;
        pixel_data[165][44] = 1;
        pixel_data[165][45] = 1;
        pixel_data[165][46] = 1;
        pixel_data[165][47] = 1;
        pixel_data[165][48] = 1;
        pixel_data[165][49] = 1;
        pixel_data[165][50] = 1;
        pixel_data[165][51] = 1;
        pixel_data[165][52] = 1;
        pixel_data[165][53] = 1;
        pixel_data[165][54] = 1;
        pixel_data[165][55] = 1;
        pixel_data[165][56] = 1;
        pixel_data[165][57] = 1;
        pixel_data[165][58] = 1;
        pixel_data[165][59] = 1;
        pixel_data[165][60] = 1;
        pixel_data[165][61] = 1;
        pixel_data[165][62] = 1;
        pixel_data[165][63] = 1;
        pixel_data[165][64] = 1;
        pixel_data[165][65] = 1;
        pixel_data[165][66] = 1;
        pixel_data[165][67] = 1;
        pixel_data[165][68] = 1;
        pixel_data[165][69] = 1;
        pixel_data[165][70] = 1;
        pixel_data[165][71] = 1;
        pixel_data[165][72] = 1;
        pixel_data[165][73] = 1;
        pixel_data[165][74] = 1;
        pixel_data[165][75] = 1;
        pixel_data[165][76] = 1;
        pixel_data[165][77] = 1;
        pixel_data[165][78] = 1;
        pixel_data[165][79] = 1;
        pixel_data[165][80] = 1;
        pixel_data[165][81] = 1;
        pixel_data[165][82] = 1;
        pixel_data[165][83] = 1;
        pixel_data[165][84] = 1;
        pixel_data[165][85] = 1;
        pixel_data[165][86] = 6;
        pixel_data[165][87] = 12;
        pixel_data[165][88] = 13;
        pixel_data[165][89] = 13;
        pixel_data[165][90] = 13;
        pixel_data[165][91] = 13;
        pixel_data[165][92] = 13;
        pixel_data[165][93] = 13;
        pixel_data[165][94] = 13;
        pixel_data[165][95] = 13;
        pixel_data[165][96] = 13;
        pixel_data[165][97] = 13;
        pixel_data[165][98] = 13;
        pixel_data[165][99] = 13;
        pixel_data[165][100] = 13;
        pixel_data[165][101] = 13;
        pixel_data[165][102] = 13;
        pixel_data[165][103] = 13;
        pixel_data[165][104] = 13;
        pixel_data[165][105] = 13;
        pixel_data[165][106] = 13;
        pixel_data[165][107] = 13;
        pixel_data[165][108] = 13;
        pixel_data[165][109] = 13;
        pixel_data[165][110] = 13;
        pixel_data[165][111] = 13;
        pixel_data[165][112] = 13;
        pixel_data[165][113] = 13;
        pixel_data[165][114] = 13;
        pixel_data[165][115] = 13;
        pixel_data[165][116] = 10;
        pixel_data[165][117] = 1;
        pixel_data[165][118] = 1;
        pixel_data[165][119] = 1;
        pixel_data[165][120] = 1;
        pixel_data[165][121] = 1;
        pixel_data[165][122] = 1;
        pixel_data[165][123] = 1;
        pixel_data[165][124] = 1;
        pixel_data[165][125] = 1;
        pixel_data[165][126] = 1;
        pixel_data[165][127] = 1;
        pixel_data[165][128] = 1;
        pixel_data[165][129] = 4;
        pixel_data[165][130] = 8;
        pixel_data[165][131] = 13;
        pixel_data[165][132] = 13;
        pixel_data[165][133] = 13;
        pixel_data[165][134] = 13;
        pixel_data[165][135] = 13;
        pixel_data[165][136] = 13;
        pixel_data[165][137] = 13;
        pixel_data[165][138] = 13;
        pixel_data[165][139] = 13;
        pixel_data[165][140] = 13;
        pixel_data[165][141] = 13;
        pixel_data[165][142] = 13;
        pixel_data[165][143] = 13;
        pixel_data[165][144] = 13;
        pixel_data[165][145] = 13;
        pixel_data[165][146] = 13;
        pixel_data[165][147] = 13;
        pixel_data[165][148] = 13;
        pixel_data[165][149] = 13;
        pixel_data[165][150] = 13;
        pixel_data[165][151] = 13;
        pixel_data[165][152] = 13;
        pixel_data[165][153] = 10;
        pixel_data[165][154] = 5;
        pixel_data[165][155] = 1;
        pixel_data[165][156] = 1;
        pixel_data[165][157] = 1;
        pixel_data[165][158] = 1;
        pixel_data[165][159] = 1;
        pixel_data[165][160] = 1;
        pixel_data[165][161] = 1;
        pixel_data[165][162] = 1;
        pixel_data[165][163] = 1;
        pixel_data[165][164] = 1;
        pixel_data[165][165] = 1;
        pixel_data[165][166] = 1;
        pixel_data[165][167] = 1;
        pixel_data[165][168] = 1;
        pixel_data[165][169] = 1;
        pixel_data[165][170] = 1;
        pixel_data[165][171] = 1;
        pixel_data[165][172] = 1;
        pixel_data[165][173] = 1;
        pixel_data[165][174] = 1;
        pixel_data[165][175] = 1;
        pixel_data[165][176] = 4;
        pixel_data[165][177] = 7;
        pixel_data[165][178] = 9;
        pixel_data[165][179] = 11;
        pixel_data[165][180] = 11;
        pixel_data[165][181] = 0;
        pixel_data[165][182] = 0;
        pixel_data[165][183] = 0;
        pixel_data[165][184] = 0;
        pixel_data[165][185] = 0;
        pixel_data[165][186] = 0;
        pixel_data[165][187] = 0;
        pixel_data[165][188] = 0;
        pixel_data[165][189] = 0;
        pixel_data[165][190] = 0;
        pixel_data[165][191] = 0;
        pixel_data[165][192] = 0;
        pixel_data[165][193] = 0;
        pixel_data[165][194] = 0;
        pixel_data[165][195] = 0;
        pixel_data[165][196] = 0;
        pixel_data[165][197] = 0;
        pixel_data[165][198] = 0;
        pixel_data[165][199] = 0; // y=165
        pixel_data[166][0] = 0;
        pixel_data[166][1] = 0;
        pixel_data[166][2] = 0;
        pixel_data[166][3] = 0;
        pixel_data[166][4] = 0;
        pixel_data[166][5] = 0;
        pixel_data[166][6] = 0;
        pixel_data[166][7] = 0;
        pixel_data[166][8] = 0;
        pixel_data[166][9] = 0;
        pixel_data[166][10] = 10;
        pixel_data[166][11] = 11;
        pixel_data[166][12] = 9;
        pixel_data[166][13] = 7;
        pixel_data[166][14] = 4;
        pixel_data[166][15] = 4;
        pixel_data[166][16] = 2;
        pixel_data[166][17] = 1;
        pixel_data[166][18] = 1;
        pixel_data[166][19] = 1;
        pixel_data[166][20] = 1;
        pixel_data[166][21] = 1;
        pixel_data[166][22] = 1;
        pixel_data[166][23] = 1;
        pixel_data[166][24] = 1;
        pixel_data[166][25] = 1;
        pixel_data[166][26] = 1;
        pixel_data[166][27] = 1;
        pixel_data[166][28] = 1;
        pixel_data[166][29] = 1;
        pixel_data[166][30] = 1;
        pixel_data[166][31] = 1;
        pixel_data[166][32] = 1;
        pixel_data[166][33] = 1;
        pixel_data[166][34] = 1;
        pixel_data[166][35] = 1;
        pixel_data[166][36] = 1;
        pixel_data[166][37] = 1;
        pixel_data[166][38] = 1;
        pixel_data[166][39] = 1;
        pixel_data[166][40] = 1;
        pixel_data[166][41] = 1;
        pixel_data[166][42] = 1;
        pixel_data[166][43] = 1;
        pixel_data[166][44] = 1;
        pixel_data[166][45] = 1;
        pixel_data[166][46] = 1;
        pixel_data[166][47] = 1;
        pixel_data[166][48] = 1;
        pixel_data[166][49] = 1;
        pixel_data[166][50] = 1;
        pixel_data[166][51] = 1;
        pixel_data[166][52] = 1;
        pixel_data[166][53] = 1;
        pixel_data[166][54] = 1;
        pixel_data[166][55] = 1;
        pixel_data[166][56] = 1;
        pixel_data[166][57] = 1;
        pixel_data[166][58] = 1;
        pixel_data[166][59] = 1;
        pixel_data[166][60] = 1;
        pixel_data[166][61] = 1;
        pixel_data[166][62] = 1;
        pixel_data[166][63] = 1;
        pixel_data[166][64] = 1;
        pixel_data[166][65] = 1;
        pixel_data[166][66] = 1;
        pixel_data[166][67] = 1;
        pixel_data[166][68] = 1;
        pixel_data[166][69] = 1;
        pixel_data[166][70] = 1;
        pixel_data[166][71] = 1;
        pixel_data[166][72] = 1;
        pixel_data[166][73] = 1;
        pixel_data[166][74] = 1;
        pixel_data[166][75] = 1;
        pixel_data[166][76] = 1;
        pixel_data[166][77] = 1;
        pixel_data[166][78] = 2;
        pixel_data[166][79] = 1;
        pixel_data[166][80] = 1;
        pixel_data[166][81] = 1;
        pixel_data[166][82] = 1;
        pixel_data[166][83] = 1;
        pixel_data[166][84] = 1;
        pixel_data[166][85] = 1;
        pixel_data[166][86] = 1;
        pixel_data[166][87] = 7;
        pixel_data[166][88] = 12;
        pixel_data[166][89] = 13;
        pixel_data[166][90] = 13;
        pixel_data[166][91] = 13;
        pixel_data[166][92] = 13;
        pixel_data[166][93] = 13;
        pixel_data[166][94] = 13;
        pixel_data[166][95] = 13;
        pixel_data[166][96] = 13;
        pixel_data[166][97] = 13;
        pixel_data[166][98] = 13;
        pixel_data[166][99] = 13;
        pixel_data[166][100] = 13;
        pixel_data[166][101] = 13;
        pixel_data[166][102] = 13;
        pixel_data[166][103] = 13;
        pixel_data[166][104] = 13;
        pixel_data[166][105] = 13;
        pixel_data[166][106] = 13;
        pixel_data[166][107] = 13;
        pixel_data[166][108] = 13;
        pixel_data[166][109] = 13;
        pixel_data[166][110] = 13;
        pixel_data[166][111] = 13;
        pixel_data[166][112] = 13;
        pixel_data[166][113] = 13;
        pixel_data[166][114] = 13;
        pixel_data[166][115] = 13;
        pixel_data[166][116] = 7;
        pixel_data[166][117] = 1;
        pixel_data[166][118] = 1;
        pixel_data[166][119] = 1;
        pixel_data[166][120] = 1;
        pixel_data[166][121] = 1;
        pixel_data[166][122] = 1;
        pixel_data[166][123] = 1;
        pixel_data[166][124] = 1;
        pixel_data[166][125] = 1;
        pixel_data[166][126] = 1;
        pixel_data[166][127] = 1;
        pixel_data[166][128] = 1;
        pixel_data[166][129] = 1;
        pixel_data[166][130] = 1;
        pixel_data[166][131] = 7;
        pixel_data[166][132] = 12;
        pixel_data[166][133] = 13;
        pixel_data[166][134] = 13;
        pixel_data[166][135] = 13;
        pixel_data[166][136] = 13;
        pixel_data[166][137] = 13;
        pixel_data[166][138] = 13;
        pixel_data[166][139] = 13;
        pixel_data[166][140] = 13;
        pixel_data[166][141] = 13;
        pixel_data[166][142] = 13;
        pixel_data[166][143] = 13;
        pixel_data[166][144] = 13;
        pixel_data[166][145] = 13;
        pixel_data[166][146] = 13;
        pixel_data[166][147] = 13;
        pixel_data[166][148] = 13;
        pixel_data[166][149] = 13;
        pixel_data[166][150] = 13;
        pixel_data[166][151] = 13;
        pixel_data[166][152] = 13;
        pixel_data[166][153] = 10;
        pixel_data[166][154] = 2;
        pixel_data[166][155] = 1;
        pixel_data[166][156] = 1;
        pixel_data[166][157] = 1;
        pixel_data[166][158] = 1;
        pixel_data[166][159] = 1;
        pixel_data[166][160] = 1;
        pixel_data[166][161] = 1;
        pixel_data[166][162] = 1;
        pixel_data[166][163] = 1;
        pixel_data[166][164] = 1;
        pixel_data[166][165] = 1;
        pixel_data[166][166] = 1;
        pixel_data[166][167] = 1;
        pixel_data[166][168] = 1;
        pixel_data[166][169] = 1;
        pixel_data[166][170] = 1;
        pixel_data[166][171] = 1;
        pixel_data[166][172] = 1;
        pixel_data[166][173] = 1;
        pixel_data[166][174] = 1;
        pixel_data[166][175] = 1;
        pixel_data[166][176] = 1;
        pixel_data[166][177] = 1;
        pixel_data[166][178] = 6;
        pixel_data[166][179] = 9;
        pixel_data[166][180] = 11;
        pixel_data[166][181] = 11;
        pixel_data[166][182] = 0;
        pixel_data[166][183] = 0;
        pixel_data[166][184] = 0;
        pixel_data[166][185] = 0;
        pixel_data[166][186] = 0;
        pixel_data[166][187] = 0;
        pixel_data[166][188] = 0;
        pixel_data[166][189] = 0;
        pixel_data[166][190] = 0;
        pixel_data[166][191] = 0;
        pixel_data[166][192] = 0;
        pixel_data[166][193] = 0;
        pixel_data[166][194] = 0;
        pixel_data[166][195] = 0;
        pixel_data[166][196] = 0;
        pixel_data[166][197] = 0;
        pixel_data[166][198] = 0;
        pixel_data[166][199] = 0; // y=166
        pixel_data[167][0] = 0;
        pixel_data[167][1] = 0;
        pixel_data[167][2] = 0;
        pixel_data[167][3] = 0;
        pixel_data[167][4] = 0;
        pixel_data[167][5] = 0;
        pixel_data[167][6] = 0;
        pixel_data[167][7] = 0;
        pixel_data[167][8] = 0;
        pixel_data[167][9] = 11;
        pixel_data[167][10] = 11;
        pixel_data[167][11] = 9;
        pixel_data[167][12] = 7;
        pixel_data[167][13] = 4;
        pixel_data[167][14] = 4;
        pixel_data[167][15] = 4;
        pixel_data[167][16] = 1;
        pixel_data[167][17] = 1;
        pixel_data[167][18] = 1;
        pixel_data[167][19] = 1;
        pixel_data[167][20] = 1;
        pixel_data[167][21] = 1;
        pixel_data[167][22] = 1;
        pixel_data[167][23] = 1;
        pixel_data[167][24] = 1;
        pixel_data[167][25] = 1;
        pixel_data[167][26] = 1;
        pixel_data[167][27] = 1;
        pixel_data[167][28] = 1;
        pixel_data[167][29] = 1;
        pixel_data[167][30] = 1;
        pixel_data[167][31] = 1;
        pixel_data[167][32] = 1;
        pixel_data[167][33] = 1;
        pixel_data[167][34] = 1;
        pixel_data[167][35] = 1;
        pixel_data[167][36] = 1;
        pixel_data[167][37] = 1;
        pixel_data[167][38] = 1;
        pixel_data[167][39] = 1;
        pixel_data[167][40] = 1;
        pixel_data[167][41] = 1;
        pixel_data[167][42] = 1;
        pixel_data[167][43] = 1;
        pixel_data[167][44] = 1;
        pixel_data[167][45] = 1;
        pixel_data[167][46] = 1;
        pixel_data[167][47] = 1;
        pixel_data[167][48] = 1;
        pixel_data[167][49] = 1;
        pixel_data[167][50] = 1;
        pixel_data[167][51] = 1;
        pixel_data[167][52] = 1;
        pixel_data[167][53] = 1;
        pixel_data[167][54] = 1;
        pixel_data[167][55] = 1;
        pixel_data[167][56] = 1;
        pixel_data[167][57] = 1;
        pixel_data[167][58] = 1;
        pixel_data[167][59] = 1;
        pixel_data[167][60] = 1;
        pixel_data[167][61] = 1;
        pixel_data[167][62] = 1;
        pixel_data[167][63] = 1;
        pixel_data[167][64] = 1;
        pixel_data[167][65] = 1;
        pixel_data[167][66] = 1;
        pixel_data[167][67] = 1;
        pixel_data[167][68] = 1;
        pixel_data[167][69] = 1;
        pixel_data[167][70] = 1;
        pixel_data[167][71] = 1;
        pixel_data[167][72] = 1;
        pixel_data[167][73] = 1;
        pixel_data[167][74] = 1;
        pixel_data[167][75] = 1;
        pixel_data[167][76] = 1;
        pixel_data[167][77] = 1;
        pixel_data[167][78] = 1;
        pixel_data[167][79] = 1;
        pixel_data[167][80] = 1;
        pixel_data[167][81] = 1;
        pixel_data[167][82] = 1;
        pixel_data[167][83] = 1;
        pixel_data[167][84] = 1;
        pixel_data[167][85] = 1;
        pixel_data[167][86] = 1;
        pixel_data[167][87] = 1;
        pixel_data[167][88] = 7;
        pixel_data[167][89] = 12;
        pixel_data[167][90] = 13;
        pixel_data[167][91] = 13;
        pixel_data[167][92] = 13;
        pixel_data[167][93] = 13;
        pixel_data[167][94] = 13;
        pixel_data[167][95] = 13;
        pixel_data[167][96] = 13;
        pixel_data[167][97] = 13;
        pixel_data[167][98] = 13;
        pixel_data[167][99] = 13;
        pixel_data[167][100] = 13;
        pixel_data[167][101] = 13;
        pixel_data[167][102] = 13;
        pixel_data[167][103] = 13;
        pixel_data[167][104] = 13;
        pixel_data[167][105] = 13;
        pixel_data[167][106] = 13;
        pixel_data[167][107] = 13;
        pixel_data[167][108] = 13;
        pixel_data[167][109] = 13;
        pixel_data[167][110] = 13;
        pixel_data[167][111] = 13;
        pixel_data[167][112] = 13;
        pixel_data[167][113] = 13;
        pixel_data[167][114] = 13;
        pixel_data[167][115] = 8;
        pixel_data[167][116] = 1;
        pixel_data[167][117] = 1;
        pixel_data[167][118] = 1;
        pixel_data[167][119] = 1;
        pixel_data[167][120] = 1;
        pixel_data[167][121] = 1;
        pixel_data[167][122] = 1;
        pixel_data[167][123] = 1;
        pixel_data[167][124] = 1;
        pixel_data[167][125] = 1;
        pixel_data[167][126] = 1;
        pixel_data[167][127] = 1;
        pixel_data[167][128] = 1;
        pixel_data[167][129] = 1;
        pixel_data[167][130] = 1;
        pixel_data[167][131] = 1;
        pixel_data[167][132] = 7;
        pixel_data[167][133] = 10;
        pixel_data[167][134] = 13;
        pixel_data[167][135] = 13;
        pixel_data[167][136] = 13;
        pixel_data[167][137] = 13;
        pixel_data[167][138] = 13;
        pixel_data[167][139] = 13;
        pixel_data[167][140] = 13;
        pixel_data[167][141] = 13;
        pixel_data[167][142] = 13;
        pixel_data[167][143] = 13;
        pixel_data[167][144] = 13;
        pixel_data[167][145] = 13;
        pixel_data[167][146] = 13;
        pixel_data[167][147] = 13;
        pixel_data[167][148] = 13;
        pixel_data[167][149] = 13;
        pixel_data[167][150] = 13;
        pixel_data[167][151] = 13;
        pixel_data[167][152] = 12;
        pixel_data[167][153] = 6;
        pixel_data[167][154] = 1;
        pixel_data[167][155] = 1;
        pixel_data[167][156] = 1;
        pixel_data[167][157] = 1;
        pixel_data[167][158] = 1;
        pixel_data[167][159] = 1;
        pixel_data[167][160] = 1;
        pixel_data[167][161] = 1;
        pixel_data[167][162] = 1;
        pixel_data[167][163] = 1;
        pixel_data[167][164] = 1;
        pixel_data[167][165] = 1;
        pixel_data[167][166] = 1;
        pixel_data[167][167] = 1;
        pixel_data[167][168] = 1;
        pixel_data[167][169] = 1;
        pixel_data[167][170] = 1;
        pixel_data[167][171] = 1;
        pixel_data[167][172] = 1;
        pixel_data[167][173] = 1;
        pixel_data[167][174] = 1;
        pixel_data[167][175] = 1;
        pixel_data[167][176] = 1;
        pixel_data[167][177] = 1;
        pixel_data[167][178] = 1;
        pixel_data[167][179] = 6;
        pixel_data[167][180] = 9;
        pixel_data[167][181] = 11;
        pixel_data[167][182] = 11;
        pixel_data[167][183] = 0;
        pixel_data[167][184] = 0;
        pixel_data[167][185] = 0;
        pixel_data[167][186] = 0;
        pixel_data[167][187] = 0;
        pixel_data[167][188] = 0;
        pixel_data[167][189] = 0;
        pixel_data[167][190] = 0;
        pixel_data[167][191] = 0;
        pixel_data[167][192] = 0;
        pixel_data[167][193] = 0;
        pixel_data[167][194] = 0;
        pixel_data[167][195] = 0;
        pixel_data[167][196] = 0;
        pixel_data[167][197] = 0;
        pixel_data[167][198] = 0;
        pixel_data[167][199] = 0; // y=167
        pixel_data[168][0] = 0;
        pixel_data[168][1] = 0;
        pixel_data[168][2] = 0;
        pixel_data[168][3] = 0;
        pixel_data[168][4] = 0;
        pixel_data[168][5] = 0;
        pixel_data[168][6] = 0;
        pixel_data[168][7] = 0;
        pixel_data[168][8] = 0;
        pixel_data[168][9] = 11;
        pixel_data[168][10] = 11;
        pixel_data[168][11] = 8;
        pixel_data[168][12] = 4;
        pixel_data[168][13] = 2;
        pixel_data[168][14] = 4;
        pixel_data[168][15] = 4;
        pixel_data[168][16] = 1;
        pixel_data[168][17] = 1;
        pixel_data[168][18] = 1;
        pixel_data[168][19] = 1;
        pixel_data[168][20] = 1;
        pixel_data[168][21] = 1;
        pixel_data[168][22] = 1;
        pixel_data[168][23] = 1;
        pixel_data[168][24] = 1;
        pixel_data[168][25] = 1;
        pixel_data[168][26] = 1;
        pixel_data[168][27] = 1;
        pixel_data[168][28] = 1;
        pixel_data[168][29] = 1;
        pixel_data[168][30] = 1;
        pixel_data[168][31] = 1;
        pixel_data[168][32] = 1;
        pixel_data[168][33] = 1;
        pixel_data[168][34] = 1;
        pixel_data[168][35] = 1;
        pixel_data[168][36] = 1;
        pixel_data[168][37] = 1;
        pixel_data[168][38] = 1;
        pixel_data[168][39] = 1;
        pixel_data[168][40] = 1;
        pixel_data[168][41] = 1;
        pixel_data[168][42] = 1;
        pixel_data[168][43] = 1;
        pixel_data[168][44] = 1;
        pixel_data[168][45] = 1;
        pixel_data[168][46] = 1;
        pixel_data[168][47] = 1;
        pixel_data[168][48] = 1;
        pixel_data[168][49] = 1;
        pixel_data[168][50] = 1;
        pixel_data[168][51] = 1;
        pixel_data[168][52] = 1;
        pixel_data[168][53] = 1;
        pixel_data[168][54] = 1;
        pixel_data[168][55] = 1;
        pixel_data[168][56] = 1;
        pixel_data[168][57] = 1;
        pixel_data[168][58] = 1;
        pixel_data[168][59] = 1;
        pixel_data[168][60] = 1;
        pixel_data[168][61] = 1;
        pixel_data[168][62] = 1;
        pixel_data[168][63] = 1;
        pixel_data[168][64] = 1;
        pixel_data[168][65] = 1;
        pixel_data[168][66] = 1;
        pixel_data[168][67] = 1;
        pixel_data[168][68] = 1;
        pixel_data[168][69] = 1;
        pixel_data[168][70] = 1;
        pixel_data[168][71] = 1;
        pixel_data[168][72] = 2;
        pixel_data[168][73] = 1;
        pixel_data[168][74] = 1;
        pixel_data[168][75] = 1;
        pixel_data[168][76] = 1;
        pixel_data[168][77] = 1;
        pixel_data[168][78] = 1;
        pixel_data[168][79] = 1;
        pixel_data[168][80] = 1;
        pixel_data[168][81] = 1;
        pixel_data[168][82] = 1;
        pixel_data[168][83] = 1;
        pixel_data[168][84] = 1;
        pixel_data[168][85] = 1;
        pixel_data[168][86] = 1;
        pixel_data[168][87] = 1;
        pixel_data[168][88] = 1;
        pixel_data[168][89] = 4;
        pixel_data[168][90] = 8;
        pixel_data[168][91] = 12;
        pixel_data[168][92] = 13;
        pixel_data[168][93] = 13;
        pixel_data[168][94] = 13;
        pixel_data[168][95] = 13;
        pixel_data[168][96] = 13;
        pixel_data[168][97] = 13;
        pixel_data[168][98] = 13;
        pixel_data[168][99] = 13;
        pixel_data[168][100] = 13;
        pixel_data[168][101] = 13;
        pixel_data[168][102] = 13;
        pixel_data[168][103] = 13;
        pixel_data[168][104] = 13;
        pixel_data[168][105] = 13;
        pixel_data[168][106] = 13;
        pixel_data[168][107] = 13;
        pixel_data[168][108] = 13;
        pixel_data[168][109] = 13;
        pixel_data[168][110] = 13;
        pixel_data[168][111] = 13;
        pixel_data[168][112] = 13;
        pixel_data[168][113] = 12;
        pixel_data[168][114] = 8;
        pixel_data[168][115] = 1;
        pixel_data[168][116] = 1;
        pixel_data[168][117] = 1;
        pixel_data[168][118] = 1;
        pixel_data[168][119] = 1;
        pixel_data[168][120] = 1;
        pixel_data[168][121] = 1;
        pixel_data[168][122] = 1;
        pixel_data[168][123] = 1;
        pixel_data[168][124] = 1;
        pixel_data[168][125] = 1;
        pixel_data[168][126] = 1;
        pixel_data[168][127] = 1;
        pixel_data[168][128] = 1;
        pixel_data[168][129] = 1;
        pixel_data[168][130] = 1;
        pixel_data[168][131] = 1;
        pixel_data[168][132] = 1;
        pixel_data[168][133] = 2;
        pixel_data[168][134] = 7;
        pixel_data[168][135] = 10;
        pixel_data[168][136] = 13;
        pixel_data[168][137] = 13;
        pixel_data[168][138] = 13;
        pixel_data[168][139] = 13;
        pixel_data[168][140] = 13;
        pixel_data[168][141] = 13;
        pixel_data[168][142] = 13;
        pixel_data[168][143] = 13;
        pixel_data[168][144] = 13;
        pixel_data[168][145] = 13;
        pixel_data[168][146] = 13;
        pixel_data[168][147] = 13;
        pixel_data[168][148] = 13;
        pixel_data[168][149] = 13;
        pixel_data[168][150] = 13;
        pixel_data[168][151] = 10;
        pixel_data[168][152] = 5;
        pixel_data[168][153] = 1;
        pixel_data[168][154] = 1;
        pixel_data[168][155] = 1;
        pixel_data[168][156] = 1;
        pixel_data[168][157] = 1;
        pixel_data[168][158] = 1;
        pixel_data[168][159] = 1;
        pixel_data[168][160] = 1;
        pixel_data[168][161] = 1;
        pixel_data[168][162] = 1;
        pixel_data[168][163] = 1;
        pixel_data[168][164] = 1;
        pixel_data[168][165] = 1;
        pixel_data[168][166] = 1;
        pixel_data[168][167] = 1;
        pixel_data[168][168] = 1;
        pixel_data[168][169] = 1;
        pixel_data[168][170] = 1;
        pixel_data[168][171] = 1;
        pixel_data[168][172] = 1;
        pixel_data[168][173] = 1;
        pixel_data[168][174] = 1;
        pixel_data[168][175] = 1;
        pixel_data[168][176] = 1;
        pixel_data[168][177] = 1;
        pixel_data[168][178] = 1;
        pixel_data[168][179] = 2;
        pixel_data[168][180] = 7;
        pixel_data[168][181] = 9;
        pixel_data[168][182] = 11;
        pixel_data[168][183] = 11;
        pixel_data[168][184] = 0;
        pixel_data[168][185] = 0;
        pixel_data[168][186] = 0;
        pixel_data[168][187] = 0;
        pixel_data[168][188] = 0;
        pixel_data[168][189] = 0;
        pixel_data[168][190] = 0;
        pixel_data[168][191] = 0;
        pixel_data[168][192] = 0;
        pixel_data[168][193] = 0;
        pixel_data[168][194] = 0;
        pixel_data[168][195] = 0;
        pixel_data[168][196] = 0;
        pixel_data[168][197] = 0;
        pixel_data[168][198] = 0;
        pixel_data[168][199] = 0; // y=168
        pixel_data[169][0] = 0;
        pixel_data[169][1] = 0;
        pixel_data[169][2] = 0;
        pixel_data[169][3] = 0;
        pixel_data[169][4] = 0;
        pixel_data[169][5] = 0;
        pixel_data[169][6] = 0;
        pixel_data[169][7] = 0;
        pixel_data[169][8] = 11;
        pixel_data[169][9] = 11;
        pixel_data[169][10] = 8;
        pixel_data[169][11] = 5;
        pixel_data[169][12] = 1;
        pixel_data[169][13] = 4;
        pixel_data[169][14] = 4;
        pixel_data[169][15] = 2;
        pixel_data[169][16] = 1;
        pixel_data[169][17] = 1;
        pixel_data[169][18] = 1;
        pixel_data[169][19] = 1;
        pixel_data[169][20] = 1;
        pixel_data[169][21] = 1;
        pixel_data[169][22] = 1;
        pixel_data[169][23] = 1;
        pixel_data[169][24] = 1;
        pixel_data[169][25] = 1;
        pixel_data[169][26] = 1;
        pixel_data[169][27] = 1;
        pixel_data[169][28] = 1;
        pixel_data[169][29] = 1;
        pixel_data[169][30] = 1;
        pixel_data[169][31] = 1;
        pixel_data[169][32] = 1;
        pixel_data[169][33] = 1;
        pixel_data[169][34] = 1;
        pixel_data[169][35] = 1;
        pixel_data[169][36] = 1;
        pixel_data[169][37] = 1;
        pixel_data[169][38] = 1;
        pixel_data[169][39] = 1;
        pixel_data[169][40] = 1;
        pixel_data[169][41] = 1;
        pixel_data[169][42] = 1;
        pixel_data[169][43] = 1;
        pixel_data[169][44] = 1;
        pixel_data[169][45] = 1;
        pixel_data[169][46] = 1;
        pixel_data[169][47] = 1;
        pixel_data[169][48] = 1;
        pixel_data[169][49] = 1;
        pixel_data[169][50] = 1;
        pixel_data[169][51] = 1;
        pixel_data[169][52] = 1;
        pixel_data[169][53] = 1;
        pixel_data[169][54] = 1;
        pixel_data[169][55] = 1;
        pixel_data[169][56] = 1;
        pixel_data[169][57] = 1;
        pixel_data[169][58] = 1;
        pixel_data[169][59] = 1;
        pixel_data[169][60] = 1;
        pixel_data[169][61] = 1;
        pixel_data[169][62] = 1;
        pixel_data[169][63] = 1;
        pixel_data[169][64] = 1;
        pixel_data[169][65] = 1;
        pixel_data[169][66] = 1;
        pixel_data[169][67] = 1;
        pixel_data[169][68] = 1;
        pixel_data[169][69] = 1;
        pixel_data[169][70] = 1;
        pixel_data[169][71] = 1;
        pixel_data[169][72] = 1;
        pixel_data[169][73] = 1;
        pixel_data[169][74] = 1;
        pixel_data[169][75] = 1;
        pixel_data[169][76] = 1;
        pixel_data[169][77] = 1;
        pixel_data[169][78] = 1;
        pixel_data[169][79] = 1;
        pixel_data[169][80] = 1;
        pixel_data[169][81] = 1;
        pixel_data[169][82] = 1;
        pixel_data[169][83] = 1;
        pixel_data[169][84] = 1;
        pixel_data[169][85] = 1;
        pixel_data[169][86] = 1;
        pixel_data[169][87] = 1;
        pixel_data[169][88] = 1;
        pixel_data[169][89] = 1;
        pixel_data[169][90] = 1;
        pixel_data[169][91] = 1;
        pixel_data[169][92] = 1;
        pixel_data[169][93] = 4;
        pixel_data[169][94] = 7;
        pixel_data[169][95] = 10;
        pixel_data[169][96] = 12;
        pixel_data[169][97] = 13;
        pixel_data[169][98] = 13;
        pixel_data[169][99] = 13;
        pixel_data[169][100] = 13;
        pixel_data[169][101] = 13;
        pixel_data[169][102] = 13;
        pixel_data[169][103] = 13;
        pixel_data[169][104] = 13;
        pixel_data[169][105] = 13;
        pixel_data[169][106] = 13;
        pixel_data[169][107] = 13;
        pixel_data[169][108] = 13;
        pixel_data[169][109] = 13;
        pixel_data[169][110] = 13;
        pixel_data[169][111] = 12;
        pixel_data[169][112] = 7;
        pixel_data[169][113] = 2;
        pixel_data[169][114] = 1;
        pixel_data[169][115] = 1;
        pixel_data[169][116] = 1;
        pixel_data[169][117] = 1;
        pixel_data[169][118] = 1;
        pixel_data[169][119] = 1;
        pixel_data[169][120] = 1;
        pixel_data[169][121] = 1;
        pixel_data[169][122] = 1;
        pixel_data[169][123] = 1;
        pixel_data[169][124] = 1;
        pixel_data[169][125] = 1;
        pixel_data[169][126] = 1;
        pixel_data[169][127] = 1;
        pixel_data[169][128] = 1;
        pixel_data[169][129] = 1;
        pixel_data[169][130] = 1;
        pixel_data[169][131] = 1;
        pixel_data[169][132] = 1;
        pixel_data[169][133] = 1;
        pixel_data[169][134] = 1;
        pixel_data[169][135] = 1;
        pixel_data[169][136] = 1;
        pixel_data[169][137] = 1;
        pixel_data[169][138] = 5;
        pixel_data[169][139] = 5;
        pixel_data[169][140] = 5;
        pixel_data[169][141] = 4;
        pixel_data[169][142] = 5;
        pixel_data[169][143] = 6;
        pixel_data[169][144] = 7;
        pixel_data[169][145] = 7;
        pixel_data[169][146] = 7;
        pixel_data[169][147] = 6;
        pixel_data[169][148] = 5;
        pixel_data[169][149] = 1;
        pixel_data[169][150] = 1;
        pixel_data[169][151] = 1;
        pixel_data[169][152] = 1;
        pixel_data[169][153] = 1;
        pixel_data[169][154] = 1;
        pixel_data[169][155] = 1;
        pixel_data[169][156] = 1;
        pixel_data[169][157] = 1;
        pixel_data[169][158] = 1;
        pixel_data[169][159] = 1;
        pixel_data[169][160] = 1;
        pixel_data[169][161] = 1;
        pixel_data[169][162] = 1;
        pixel_data[169][163] = 1;
        pixel_data[169][164] = 1;
        pixel_data[169][165] = 1;
        pixel_data[169][166] = 1;
        pixel_data[169][167] = 1;
        pixel_data[169][168] = 1;
        pixel_data[169][169] = 1;
        pixel_data[169][170] = 1;
        pixel_data[169][171] = 1;
        pixel_data[169][172] = 1;
        pixel_data[169][173] = 1;
        pixel_data[169][174] = 1;
        pixel_data[169][175] = 1;
        pixel_data[169][176] = 1;
        pixel_data[169][177] = 1;
        pixel_data[169][178] = 1;
        pixel_data[169][179] = 1;
        pixel_data[169][180] = 2;
        pixel_data[169][181] = 7;
        pixel_data[169][182] = 9;
        pixel_data[169][183] = 11;
        pixel_data[169][184] = 11;
        pixel_data[169][185] = 0;
        pixel_data[169][186] = 0;
        pixel_data[169][187] = 0;
        pixel_data[169][188] = 0;
        pixel_data[169][189] = 0;
        pixel_data[169][190] = 0;
        pixel_data[169][191] = 0;
        pixel_data[169][192] = 0;
        pixel_data[169][193] = 0;
        pixel_data[169][194] = 0;
        pixel_data[169][195] = 0;
        pixel_data[169][196] = 0;
        pixel_data[169][197] = 0;
        pixel_data[169][198] = 0;
        pixel_data[169][199] = 0; // y=169
        pixel_data[170][0] = 0;
        pixel_data[170][1] = 0;
        pixel_data[170][2] = 0;
        pixel_data[170][3] = 0;
        pixel_data[170][4] = 0;
        pixel_data[170][5] = 0;
        pixel_data[170][6] = 0;
        pixel_data[170][7] = 11;
        pixel_data[170][8] = 11;
        pixel_data[170][9] = 9;
        pixel_data[170][10] = 6;
        pixel_data[170][11] = 1;
        pixel_data[170][12] = 1;
        pixel_data[170][13] = 4;
        pixel_data[170][14] = 4;
        pixel_data[170][15] = 2;
        pixel_data[170][16] = 1;
        pixel_data[170][17] = 1;
        pixel_data[170][18] = 1;
        pixel_data[170][19] = 1;
        pixel_data[170][20] = 1;
        pixel_data[170][21] = 1;
        pixel_data[170][22] = 1;
        pixel_data[170][23] = 1;
        pixel_data[170][24] = 1;
        pixel_data[170][25] = 1;
        pixel_data[170][26] = 1;
        pixel_data[170][27] = 1;
        pixel_data[170][28] = 1;
        pixel_data[170][29] = 1;
        pixel_data[170][30] = 1;
        pixel_data[170][31] = 1;
        pixel_data[170][32] = 1;
        pixel_data[170][33] = 1;
        pixel_data[170][34] = 1;
        pixel_data[170][35] = 1;
        pixel_data[170][36] = 1;
        pixel_data[170][37] = 1;
        pixel_data[170][38] = 1;
        pixel_data[170][39] = 1;
        pixel_data[170][40] = 1;
        pixel_data[170][41] = 1;
        pixel_data[170][42] = 1;
        pixel_data[170][43] = 1;
        pixel_data[170][44] = 1;
        pixel_data[170][45] = 1;
        pixel_data[170][46] = 1;
        pixel_data[170][47] = 1;
        pixel_data[170][48] = 1;
        pixel_data[170][49] = 1;
        pixel_data[170][50] = 1;
        pixel_data[170][51] = 1;
        pixel_data[170][52] = 1;
        pixel_data[170][53] = 1;
        pixel_data[170][54] = 1;
        pixel_data[170][55] = 1;
        pixel_data[170][56] = 1;
        pixel_data[170][57] = 1;
        pixel_data[170][58] = 1;
        pixel_data[170][59] = 1;
        pixel_data[170][60] = 1;
        pixel_data[170][61] = 1;
        pixel_data[170][62] = 1;
        pixel_data[170][63] = 1;
        pixel_data[170][64] = 1;
        pixel_data[170][65] = 1;
        pixel_data[170][66] = 1;
        pixel_data[170][67] = 1;
        pixel_data[170][68] = 1;
        pixel_data[170][69] = 1;
        pixel_data[170][70] = 1;
        pixel_data[170][71] = 1;
        pixel_data[170][72] = 1;
        pixel_data[170][73] = 1;
        pixel_data[170][74] = 1;
        pixel_data[170][75] = 1;
        pixel_data[170][76] = 1;
        pixel_data[170][77] = 1;
        pixel_data[170][78] = 1;
        pixel_data[170][79] = 1;
        pixel_data[170][80] = 1;
        pixel_data[170][81] = 1;
        pixel_data[170][82] = 1;
        pixel_data[170][83] = 1;
        pixel_data[170][84] = 1;
        pixel_data[170][85] = 1;
        pixel_data[170][86] = 1;
        pixel_data[170][87] = 1;
        pixel_data[170][88] = 1;
        pixel_data[170][89] = 1;
        pixel_data[170][90] = 1;
        pixel_data[170][91] = 1;
        pixel_data[170][92] = 1;
        pixel_data[170][93] = 1;
        pixel_data[170][94] = 1;
        pixel_data[170][95] = 1;
        pixel_data[170][96] = 1;
        pixel_data[170][97] = 1;
        pixel_data[170][98] = 4;
        pixel_data[170][99] = 5;
        pixel_data[170][100] = 6;
        pixel_data[170][101] = 7;
        pixel_data[170][102] = 8;
        pixel_data[170][103] = 9;
        pixel_data[170][104] = 10;
        pixel_data[170][105] = 10;
        pixel_data[170][106] = 10;
        pixel_data[170][107] = 9;
        pixel_data[170][108] = 8;
        pixel_data[170][109] = 6;
        pixel_data[170][110] = 2;
        pixel_data[170][111] = 1;
        pixel_data[170][112] = 1;
        pixel_data[170][113] = 1;
        pixel_data[170][114] = 1;
        pixel_data[170][115] = 1;
        pixel_data[170][116] = 1;
        pixel_data[170][117] = 1;
        pixel_data[170][118] = 1;
        pixel_data[170][119] = 1;
        pixel_data[170][120] = 1;
        pixel_data[170][121] = 1;
        pixel_data[170][122] = 1;
        pixel_data[170][123] = 1;
        pixel_data[170][124] = 1;
        pixel_data[170][125] = 1;
        pixel_data[170][126] = 1;
        pixel_data[170][127] = 1;
        pixel_data[170][128] = 1;
        pixel_data[170][129] = 1;
        pixel_data[170][130] = 1;
        pixel_data[170][131] = 1;
        pixel_data[170][132] = 1;
        pixel_data[170][133] = 1;
        pixel_data[170][134] = 1;
        pixel_data[170][135] = 1;
        pixel_data[170][136] = 1;
        pixel_data[170][137] = 1;
        pixel_data[170][138] = 1;
        pixel_data[170][139] = 1;
        pixel_data[170][140] = 1;
        pixel_data[170][141] = 1;
        pixel_data[170][142] = 1;
        pixel_data[170][143] = 1;
        pixel_data[170][144] = 1;
        pixel_data[170][145] = 1;
        pixel_data[170][146] = 1;
        pixel_data[170][147] = 1;
        pixel_data[170][148] = 1;
        pixel_data[170][149] = 1;
        pixel_data[170][150] = 1;
        pixel_data[170][151] = 1;
        pixel_data[170][152] = 1;
        pixel_data[170][153] = 1;
        pixel_data[170][154] = 1;
        pixel_data[170][155] = 1;
        pixel_data[170][156] = 1;
        pixel_data[170][157] = 1;
        pixel_data[170][158] = 1;
        pixel_data[170][159] = 1;
        pixel_data[170][160] = 1;
        pixel_data[170][161] = 1;
        pixel_data[170][162] = 1;
        pixel_data[170][163] = 1;
        pixel_data[170][164] = 1;
        pixel_data[170][165] = 1;
        pixel_data[170][166] = 1;
        pixel_data[170][167] = 1;
        pixel_data[170][168] = 1;
        pixel_data[170][169] = 1;
        pixel_data[170][170] = 1;
        pixel_data[170][171] = 1;
        pixel_data[170][172] = 1;
        pixel_data[170][173] = 1;
        pixel_data[170][174] = 1;
        pixel_data[170][175] = 1;
        pixel_data[170][176] = 1;
        pixel_data[170][177] = 1;
        pixel_data[170][178] = 1;
        pixel_data[170][179] = 1;
        pixel_data[170][180] = 1;
        pixel_data[170][181] = 5;
        pixel_data[170][182] = 8;
        pixel_data[170][183] = 11;
        pixel_data[170][184] = 11;
        pixel_data[170][185] = 0;
        pixel_data[170][186] = 0;
        pixel_data[170][187] = 0;
        pixel_data[170][188] = 0;
        pixel_data[170][189] = 0;
        pixel_data[170][190] = 0;
        pixel_data[170][191] = 0;
        pixel_data[170][192] = 0;
        pixel_data[170][193] = 0;
        pixel_data[170][194] = 0;
        pixel_data[170][195] = 0;
        pixel_data[170][196] = 0;
        pixel_data[170][197] = 0;
        pixel_data[170][198] = 0;
        pixel_data[170][199] = 0; // y=170
        pixel_data[171][0] = 0;
        pixel_data[171][1] = 0;
        pixel_data[171][2] = 0;
        pixel_data[171][3] = 0;
        pixel_data[171][4] = 0;
        pixel_data[171][5] = 0;
        pixel_data[171][6] = 0;
        pixel_data[171][7] = 11;
        pixel_data[171][8] = 11;
        pixel_data[171][9] = 8;
        pixel_data[171][10] = 4;
        pixel_data[171][11] = 1;
        pixel_data[171][12] = 1;
        pixel_data[171][13] = 4;
        pixel_data[171][14] = 4;
        pixel_data[171][15] = 2;
        pixel_data[171][16] = 1;
        pixel_data[171][17] = 1;
        pixel_data[171][18] = 1;
        pixel_data[171][19] = 1;
        pixel_data[171][20] = 1;
        pixel_data[171][21] = 1;
        pixel_data[171][22] = 1;
        pixel_data[171][23] = 1;
        pixel_data[171][24] = 1;
        pixel_data[171][25] = 1;
        pixel_data[171][26] = 1;
        pixel_data[171][27] = 1;
        pixel_data[171][28] = 1;
        pixel_data[171][29] = 1;
        pixel_data[171][30] = 1;
        pixel_data[171][31] = 1;
        pixel_data[171][32] = 1;
        pixel_data[171][33] = 1;
        pixel_data[171][34] = 1;
        pixel_data[171][35] = 1;
        pixel_data[171][36] = 1;
        pixel_data[171][37] = 1;
        pixel_data[171][38] = 1;
        pixel_data[171][39] = 1;
        pixel_data[171][40] = 1;
        pixel_data[171][41] = 1;
        pixel_data[171][42] = 1;
        pixel_data[171][43] = 1;
        pixel_data[171][44] = 1;
        pixel_data[171][45] = 1;
        pixel_data[171][46] = 1;
        pixel_data[171][47] = 1;
        pixel_data[171][48] = 1;
        pixel_data[171][49] = 1;
        pixel_data[171][50] = 1;
        pixel_data[171][51] = 1;
        pixel_data[171][52] = 1;
        pixel_data[171][53] = 1;
        pixel_data[171][54] = 1;
        pixel_data[171][55] = 1;
        pixel_data[171][56] = 1;
        pixel_data[171][57] = 1;
        pixel_data[171][58] = 1;
        pixel_data[171][59] = 1;
        pixel_data[171][60] = 1;
        pixel_data[171][61] = 1;
        pixel_data[171][62] = 1;
        pixel_data[171][63] = 1;
        pixel_data[171][64] = 1;
        pixel_data[171][65] = 1;
        pixel_data[171][66] = 1;
        pixel_data[171][67] = 1;
        pixel_data[171][68] = 1;
        pixel_data[171][69] = 1;
        pixel_data[171][70] = 1;
        pixel_data[171][71] = 1;
        pixel_data[171][72] = 1;
        pixel_data[171][73] = 1;
        pixel_data[171][74] = 1;
        pixel_data[171][75] = 1;
        pixel_data[171][76] = 1;
        pixel_data[171][77] = 1;
        pixel_data[171][78] = 1;
        pixel_data[171][79] = 1;
        pixel_data[171][80] = 1;
        pixel_data[171][81] = 1;
        pixel_data[171][82] = 1;
        pixel_data[171][83] = 1;
        pixel_data[171][84] = 1;
        pixel_data[171][85] = 1;
        pixel_data[171][86] = 1;
        pixel_data[171][87] = 1;
        pixel_data[171][88] = 1;
        pixel_data[171][89] = 1;
        pixel_data[171][90] = 1;
        pixel_data[171][91] = 1;
        pixel_data[171][92] = 1;
        pixel_data[171][93] = 1;
        pixel_data[171][94] = 1;
        pixel_data[171][95] = 1;
        pixel_data[171][96] = 1;
        pixel_data[171][97] = 1;
        pixel_data[171][98] = 1;
        pixel_data[171][99] = 1;
        pixel_data[171][100] = 1;
        pixel_data[171][101] = 1;
        pixel_data[171][102] = 1;
        pixel_data[171][103] = 1;
        pixel_data[171][104] = 1;
        pixel_data[171][105] = 1;
        pixel_data[171][106] = 1;
        pixel_data[171][107] = 1;
        pixel_data[171][108] = 1;
        pixel_data[171][109] = 1;
        pixel_data[171][110] = 1;
        pixel_data[171][111] = 1;
        pixel_data[171][112] = 1;
        pixel_data[171][113] = 1;
        pixel_data[171][114] = 1;
        pixel_data[171][115] = 1;
        pixel_data[171][116] = 1;
        pixel_data[171][117] = 1;
        pixel_data[171][118] = 1;
        pixel_data[171][119] = 1;
        pixel_data[171][120] = 1;
        pixel_data[171][121] = 1;
        pixel_data[171][122] = 1;
        pixel_data[171][123] = 1;
        pixel_data[171][124] = 1;
        pixel_data[171][125] = 1;
        pixel_data[171][126] = 1;
        pixel_data[171][127] = 1;
        pixel_data[171][128] = 1;
        pixel_data[171][129] = 1;
        pixel_data[171][130] = 1;
        pixel_data[171][131] = 1;
        pixel_data[171][132] = 1;
        pixel_data[171][133] = 1;
        pixel_data[171][134] = 1;
        pixel_data[171][135] = 1;
        pixel_data[171][136] = 1;
        pixel_data[171][137] = 1;
        pixel_data[171][138] = 1;
        pixel_data[171][139] = 1;
        pixel_data[171][140] = 1;
        pixel_data[171][141] = 1;
        pixel_data[171][142] = 1;
        pixel_data[171][143] = 1;
        pixel_data[171][144] = 1;
        pixel_data[171][145] = 1;
        pixel_data[171][146] = 1;
        pixel_data[171][147] = 1;
        pixel_data[171][148] = 1;
        pixel_data[171][149] = 1;
        pixel_data[171][150] = 1;
        pixel_data[171][151] = 1;
        pixel_data[171][152] = 1;
        pixel_data[171][153] = 1;
        pixel_data[171][154] = 1;
        pixel_data[171][155] = 1;
        pixel_data[171][156] = 1;
        pixel_data[171][157] = 1;
        pixel_data[171][158] = 1;
        pixel_data[171][159] = 1;
        pixel_data[171][160] = 1;
        pixel_data[171][161] = 1;
        pixel_data[171][162] = 1;
        pixel_data[171][163] = 1;
        pixel_data[171][164] = 1;
        pixel_data[171][165] = 1;
        pixel_data[171][166] = 1;
        pixel_data[171][167] = 1;
        pixel_data[171][168] = 1;
        pixel_data[171][169] = 1;
        pixel_data[171][170] = 1;
        pixel_data[171][171] = 1;
        pixel_data[171][172] = 1;
        pixel_data[171][173] = 1;
        pixel_data[171][174] = 1;
        pixel_data[171][175] = 1;
        pixel_data[171][176] = 1;
        pixel_data[171][177] = 1;
        pixel_data[171][178] = 1;
        pixel_data[171][179] = 1;
        pixel_data[171][180] = 1;
        pixel_data[171][181] = 1;
        pixel_data[171][182] = 7;
        pixel_data[171][183] = 9;
        pixel_data[171][184] = 11;
        pixel_data[171][185] = 10;
        pixel_data[171][186] = 0;
        pixel_data[171][187] = 0;
        pixel_data[171][188] = 0;
        pixel_data[171][189] = 0;
        pixel_data[171][190] = 0;
        pixel_data[171][191] = 0;
        pixel_data[171][192] = 0;
        pixel_data[171][193] = 0;
        pixel_data[171][194] = 0;
        pixel_data[171][195] = 0;
        pixel_data[171][196] = 0;
        pixel_data[171][197] = 0;
        pixel_data[171][198] = 0;
        pixel_data[171][199] = 0; // y=171
        pixel_data[172][0] = 0;
        pixel_data[172][1] = 0;
        pixel_data[172][2] = 0;
        pixel_data[172][3] = 0;
        pixel_data[172][4] = 0;
        pixel_data[172][5] = 0;
        pixel_data[172][6] = 11;
        pixel_data[172][7] = 11;
        pixel_data[172][8] = 8;
        pixel_data[172][9] = 6;
        pixel_data[172][10] = 1;
        pixel_data[172][11] = 1;
        pixel_data[172][12] = 2;
        pixel_data[172][13] = 4;
        pixel_data[172][14] = 4;
        pixel_data[172][15] = 1;
        pixel_data[172][16] = 1;
        pixel_data[172][17] = 1;
        pixel_data[172][18] = 1;
        pixel_data[172][19] = 1;
        pixel_data[172][20] = 1;
        pixel_data[172][21] = 1;
        pixel_data[172][22] = 1;
        pixel_data[172][23] = 1;
        pixel_data[172][24] = 1;
        pixel_data[172][25] = 1;
        pixel_data[172][26] = 1;
        pixel_data[172][27] = 1;
        pixel_data[172][28] = 1;
        pixel_data[172][29] = 1;
        pixel_data[172][30] = 1;
        pixel_data[172][31] = 1;
        pixel_data[172][32] = 1;
        pixel_data[172][33] = 1;
        pixel_data[172][34] = 1;
        pixel_data[172][35] = 1;
        pixel_data[172][36] = 1;
        pixel_data[172][37] = 1;
        pixel_data[172][38] = 1;
        pixel_data[172][39] = 1;
        pixel_data[172][40] = 1;
        pixel_data[172][41] = 1;
        pixel_data[172][42] = 1;
        pixel_data[172][43] = 1;
        pixel_data[172][44] = 1;
        pixel_data[172][45] = 1;
        pixel_data[172][46] = 1;
        pixel_data[172][47] = 1;
        pixel_data[172][48] = 1;
        pixel_data[172][49] = 1;
        pixel_data[172][50] = 1;
        pixel_data[172][51] = 1;
        pixel_data[172][52] = 1;
        pixel_data[172][53] = 1;
        pixel_data[172][54] = 1;
        pixel_data[172][55] = 1;
        pixel_data[172][56] = 1;
        pixel_data[172][57] = 1;
        pixel_data[172][58] = 1;
        pixel_data[172][59] = 1;
        pixel_data[172][60] = 1;
        pixel_data[172][61] = 1;
        pixel_data[172][62] = 1;
        pixel_data[172][63] = 1;
        pixel_data[172][64] = 1;
        pixel_data[172][65] = 1;
        pixel_data[172][66] = 1;
        pixel_data[172][67] = 1;
        pixel_data[172][68] = 1;
        pixel_data[172][69] = 1;
        pixel_data[172][70] = 1;
        pixel_data[172][71] = 1;
        pixel_data[172][72] = 1;
        pixel_data[172][73] = 1;
        pixel_data[172][74] = 1;
        pixel_data[172][75] = 1;
        pixel_data[172][76] = 1;
        pixel_data[172][77] = 1;
        pixel_data[172][78] = 1;
        pixel_data[172][79] = 1;
        pixel_data[172][80] = 1;
        pixel_data[172][81] = 1;
        pixel_data[172][82] = 1;
        pixel_data[172][83] = 1;
        pixel_data[172][84] = 1;
        pixel_data[172][85] = 1;
        pixel_data[172][86] = 1;
        pixel_data[172][87] = 1;
        pixel_data[172][88] = 1;
        pixel_data[172][89] = 1;
        pixel_data[172][90] = 1;
        pixel_data[172][91] = 1;
        pixel_data[172][92] = 1;
        pixel_data[172][93] = 1;
        pixel_data[172][94] = 1;
        pixel_data[172][95] = 1;
        pixel_data[172][96] = 1;
        pixel_data[172][97] = 1;
        pixel_data[172][98] = 1;
        pixel_data[172][99] = 1;
        pixel_data[172][100] = 1;
        pixel_data[172][101] = 1;
        pixel_data[172][102] = 1;
        pixel_data[172][103] = 1;
        pixel_data[172][104] = 1;
        pixel_data[172][105] = 1;
        pixel_data[172][106] = 1;
        pixel_data[172][107] = 1;
        pixel_data[172][108] = 1;
        pixel_data[172][109] = 1;
        pixel_data[172][110] = 1;
        pixel_data[172][111] = 1;
        pixel_data[172][112] = 1;
        pixel_data[172][113] = 1;
        pixel_data[172][114] = 1;
        pixel_data[172][115] = 1;
        pixel_data[172][116] = 1;
        pixel_data[172][117] = 1;
        pixel_data[172][118] = 1;
        pixel_data[172][119] = 1;
        pixel_data[172][120] = 1;
        pixel_data[172][121] = 1;
        pixel_data[172][122] = 1;
        pixel_data[172][123] = 1;
        pixel_data[172][124] = 1;
        pixel_data[172][125] = 1;
        pixel_data[172][126] = 1;
        pixel_data[172][127] = 1;
        pixel_data[172][128] = 1;
        pixel_data[172][129] = 1;
        pixel_data[172][130] = 1;
        pixel_data[172][131] = 1;
        pixel_data[172][132] = 1;
        pixel_data[172][133] = 1;
        pixel_data[172][134] = 1;
        pixel_data[172][135] = 1;
        pixel_data[172][136] = 1;
        pixel_data[172][137] = 1;
        pixel_data[172][138] = 1;
        pixel_data[172][139] = 1;
        pixel_data[172][140] = 1;
        pixel_data[172][141] = 1;
        pixel_data[172][142] = 1;
        pixel_data[172][143] = 1;
        pixel_data[172][144] = 1;
        pixel_data[172][145] = 1;
        pixel_data[172][146] = 1;
        pixel_data[172][147] = 1;
        pixel_data[172][148] = 1;
        pixel_data[172][149] = 1;
        pixel_data[172][150] = 1;
        pixel_data[172][151] = 1;
        pixel_data[172][152] = 1;
        pixel_data[172][153] = 1;
        pixel_data[172][154] = 1;
        pixel_data[172][155] = 1;
        pixel_data[172][156] = 1;
        pixel_data[172][157] = 1;
        pixel_data[172][158] = 1;
        pixel_data[172][159] = 1;
        pixel_data[172][160] = 1;
        pixel_data[172][161] = 1;
        pixel_data[172][162] = 1;
        pixel_data[172][163] = 1;
        pixel_data[172][164] = 1;
        pixel_data[172][165] = 1;
        pixel_data[172][166] = 1;
        pixel_data[172][167] = 1;
        pixel_data[172][168] = 1;
        pixel_data[172][169] = 1;
        pixel_data[172][170] = 1;
        pixel_data[172][171] = 1;
        pixel_data[172][172] = 1;
        pixel_data[172][173] = 1;
        pixel_data[172][174] = 1;
        pixel_data[172][175] = 1;
        pixel_data[172][176] = 1;
        pixel_data[172][177] = 1;
        pixel_data[172][178] = 1;
        pixel_data[172][179] = 1;
        pixel_data[172][180] = 1;
        pixel_data[172][181] = 1;
        pixel_data[172][182] = 2;
        pixel_data[172][183] = 7;
        pixel_data[172][184] = 9;
        pixel_data[172][185] = 11;
        pixel_data[172][186] = 11;
        pixel_data[172][187] = 0;
        pixel_data[172][188] = 0;
        pixel_data[172][189] = 0;
        pixel_data[172][190] = 0;
        pixel_data[172][191] = 0;
        pixel_data[172][192] = 0;
        pixel_data[172][193] = 0;
        pixel_data[172][194] = 0;
        pixel_data[172][195] = 0;
        pixel_data[172][196] = 0;
        pixel_data[172][197] = 0;
        pixel_data[172][198] = 0;
        pixel_data[172][199] = 0; // y=172
        pixel_data[173][0] = 0;
        pixel_data[173][1] = 0;
        pixel_data[173][2] = 0;
        pixel_data[173][3] = 0;
        pixel_data[173][4] = 0;
        pixel_data[173][5] = 13;
        pixel_data[173][6] = 11;
        pixel_data[173][7] = 11;
        pixel_data[173][8] = 7;
        pixel_data[173][9] = 1;
        pixel_data[173][10] = 1;
        pixel_data[173][11] = 1;
        pixel_data[173][12] = 2;
        pixel_data[173][13] = 4;
        pixel_data[173][14] = 4;
        pixel_data[173][15] = 1;
        pixel_data[173][16] = 1;
        pixel_data[173][17] = 1;
        pixel_data[173][18] = 1;
        pixel_data[173][19] = 1;
        pixel_data[173][20] = 1;
        pixel_data[173][21] = 1;
        pixel_data[173][22] = 1;
        pixel_data[173][23] = 1;
        pixel_data[173][24] = 1;
        pixel_data[173][25] = 1;
        pixel_data[173][26] = 1;
        pixel_data[173][27] = 1;
        pixel_data[173][28] = 1;
        pixel_data[173][29] = 1;
        pixel_data[173][30] = 1;
        pixel_data[173][31] = 1;
        pixel_data[173][32] = 1;
        pixel_data[173][33] = 1;
        pixel_data[173][34] = 1;
        pixel_data[173][35] = 1;
        pixel_data[173][36] = 1;
        pixel_data[173][37] = 1;
        pixel_data[173][38] = 1;
        pixel_data[173][39] = 1;
        pixel_data[173][40] = 1;
        pixel_data[173][41] = 1;
        pixel_data[173][42] = 1;
        pixel_data[173][43] = 1;
        pixel_data[173][44] = 1;
        pixel_data[173][45] = 1;
        pixel_data[173][46] = 1;
        pixel_data[173][47] = 1;
        pixel_data[173][48] = 1;
        pixel_data[173][49] = 1;
        pixel_data[173][50] = 1;
        pixel_data[173][51] = 1;
        pixel_data[173][52] = 1;
        pixel_data[173][53] = 1;
        pixel_data[173][54] = 1;
        pixel_data[173][55] = 1;
        pixel_data[173][56] = 1;
        pixel_data[173][57] = 1;
        pixel_data[173][58] = 1;
        pixel_data[173][59] = 1;
        pixel_data[173][60] = 1;
        pixel_data[173][61] = 1;
        pixel_data[173][62] = 1;
        pixel_data[173][63] = 1;
        pixel_data[173][64] = 1;
        pixel_data[173][65] = 1;
        pixel_data[173][66] = 1;
        pixel_data[173][67] = 1;
        pixel_data[173][68] = 1;
        pixel_data[173][69] = 1;
        pixel_data[173][70] = 1;
        pixel_data[173][71] = 1;
        pixel_data[173][72] = 1;
        pixel_data[173][73] = 1;
        pixel_data[173][74] = 1;
        pixel_data[173][75] = 1;
        pixel_data[173][76] = 1;
        pixel_data[173][77] = 1;
        pixel_data[173][78] = 1;
        pixel_data[173][79] = 1;
        pixel_data[173][80] = 1;
        pixel_data[173][81] = 1;
        pixel_data[173][82] = 1;
        pixel_data[173][83] = 1;
        pixel_data[173][84] = 1;
        pixel_data[173][85] = 1;
        pixel_data[173][86] = 1;
        pixel_data[173][87] = 1;
        pixel_data[173][88] = 1;
        pixel_data[173][89] = 1;
        pixel_data[173][90] = 1;
        pixel_data[173][91] = 1;
        pixel_data[173][92] = 1;
        pixel_data[173][93] = 1;
        pixel_data[173][94] = 1;
        pixel_data[173][95] = 1;
        pixel_data[173][96] = 1;
        pixel_data[173][97] = 1;
        pixel_data[173][98] = 1;
        pixel_data[173][99] = 1;
        pixel_data[173][100] = 1;
        pixel_data[173][101] = 1;
        pixel_data[173][102] = 1;
        pixel_data[173][103] = 1;
        pixel_data[173][104] = 1;
        pixel_data[173][105] = 1;
        pixel_data[173][106] = 1;
        pixel_data[173][107] = 1;
        pixel_data[173][108] = 1;
        pixel_data[173][109] = 1;
        pixel_data[173][110] = 1;
        pixel_data[173][111] = 1;
        pixel_data[173][112] = 1;
        pixel_data[173][113] = 1;
        pixel_data[173][114] = 1;
        pixel_data[173][115] = 1;
        pixel_data[173][116] = 1;
        pixel_data[173][117] = 1;
        pixel_data[173][118] = 1;
        pixel_data[173][119] = 1;
        pixel_data[173][120] = 1;
        pixel_data[173][121] = 1;
        pixel_data[173][122] = 1;
        pixel_data[173][123] = 6;
        pixel_data[173][124] = 9;
        pixel_data[173][125] = 10;
        pixel_data[173][126] = 8;
        pixel_data[173][127] = 5;
        pixel_data[173][128] = 1;
        pixel_data[173][129] = 1;
        pixel_data[173][130] = 1;
        pixel_data[173][131] = 1;
        pixel_data[173][132] = 1;
        pixel_data[173][133] = 1;
        pixel_data[173][134] = 1;
        pixel_data[173][135] = 1;
        pixel_data[173][136] = 1;
        pixel_data[173][137] = 1;
        pixel_data[173][138] = 1;
        pixel_data[173][139] = 1;
        pixel_data[173][140] = 1;
        pixel_data[173][141] = 1;
        pixel_data[173][142] = 1;
        pixel_data[173][143] = 1;
        pixel_data[173][144] = 1;
        pixel_data[173][145] = 1;
        pixel_data[173][146] = 1;
        pixel_data[173][147] = 1;
        pixel_data[173][148] = 1;
        pixel_data[173][149] = 1;
        pixel_data[173][150] = 1;
        pixel_data[173][151] = 1;
        pixel_data[173][152] = 1;
        pixel_data[173][153] = 1;
        pixel_data[173][154] = 1;
        pixel_data[173][155] = 1;
        pixel_data[173][156] = 1;
        pixel_data[173][157] = 1;
        pixel_data[173][158] = 1;
        pixel_data[173][159] = 1;
        pixel_data[173][160] = 1;
        pixel_data[173][161] = 1;
        pixel_data[173][162] = 1;
        pixel_data[173][163] = 1;
        pixel_data[173][164] = 1;
        pixel_data[173][165] = 1;
        pixel_data[173][166] = 1;
        pixel_data[173][167] = 1;
        pixel_data[173][168] = 1;
        pixel_data[173][169] = 1;
        pixel_data[173][170] = 1;
        pixel_data[173][171] = 1;
        pixel_data[173][172] = 1;
        pixel_data[173][173] = 1;
        pixel_data[173][174] = 1;
        pixel_data[173][175] = 1;
        pixel_data[173][176] = 1;
        pixel_data[173][177] = 1;
        pixel_data[173][178] = 1;
        pixel_data[173][179] = 1;
        pixel_data[173][180] = 1;
        pixel_data[173][181] = 1;
        pixel_data[173][182] = 1;
        pixel_data[173][183] = 5;
        pixel_data[173][184] = 8;
        pixel_data[173][185] = 11;
        pixel_data[173][186] = 11;
        pixel_data[173][187] = 0;
        pixel_data[173][188] = 0;
        pixel_data[173][189] = 0;
        pixel_data[173][190] = 0;
        pixel_data[173][191] = 0;
        pixel_data[173][192] = 0;
        pixel_data[173][193] = 0;
        pixel_data[173][194] = 0;
        pixel_data[173][195] = 0;
        pixel_data[173][196] = 0;
        pixel_data[173][197] = 0;
        pixel_data[173][198] = 0;
        pixel_data[173][199] = 0; // y=173
        pixel_data[174][0] = 0;
        pixel_data[174][1] = 0;
        pixel_data[174][2] = 0;
        pixel_data[174][3] = 0;
        pixel_data[174][4] = 0;
        pixel_data[174][5] = 11;
        pixel_data[174][6] = 11;
        pixel_data[174][7] = 9;
        pixel_data[174][8] = 6;
        pixel_data[174][9] = 1;
        pixel_data[174][10] = 1;
        pixel_data[174][11] = 1;
        pixel_data[174][12] = 2;
        pixel_data[174][13] = 4;
        pixel_data[174][14] = 4;
        pixel_data[174][15] = 1;
        pixel_data[174][16] = 1;
        pixel_data[174][17] = 1;
        pixel_data[174][18] = 1;
        pixel_data[174][19] = 1;
        pixel_data[174][20] = 1;
        pixel_data[174][21] = 1;
        pixel_data[174][22] = 1;
        pixel_data[174][23] = 1;
        pixel_data[174][24] = 1;
        pixel_data[174][25] = 1;
        pixel_data[174][26] = 1;
        pixel_data[174][27] = 1;
        pixel_data[174][28] = 1;
        pixel_data[174][29] = 1;
        pixel_data[174][30] = 1;
        pixel_data[174][31] = 1;
        pixel_data[174][32] = 1;
        pixel_data[174][33] = 1;
        pixel_data[174][34] = 1;
        pixel_data[174][35] = 1;
        pixel_data[174][36] = 1;
        pixel_data[174][37] = 1;
        pixel_data[174][38] = 1;
        pixel_data[174][39] = 1;
        pixel_data[174][40] = 1;
        pixel_data[174][41] = 1;
        pixel_data[174][42] = 1;
        pixel_data[174][43] = 1;
        pixel_data[174][44] = 1;
        pixel_data[174][45] = 1;
        pixel_data[174][46] = 1;
        pixel_data[174][47] = 1;
        pixel_data[174][48] = 1;
        pixel_data[174][49] = 1;
        pixel_data[174][50] = 1;
        pixel_data[174][51] = 1;
        pixel_data[174][52] = 1;
        pixel_data[174][53] = 1;
        pixel_data[174][54] = 1;
        pixel_data[174][55] = 1;
        pixel_data[174][56] = 1;
        pixel_data[174][57] = 1;
        pixel_data[174][58] = 1;
        pixel_data[174][59] = 1;
        pixel_data[174][60] = 1;
        pixel_data[174][61] = 1;
        pixel_data[174][62] = 1;
        pixel_data[174][63] = 1;
        pixel_data[174][64] = 1;
        pixel_data[174][65] = 1;
        pixel_data[174][66] = 1;
        pixel_data[174][67] = 1;
        pixel_data[174][68] = 1;
        pixel_data[174][69] = 1;
        pixel_data[174][70] = 1;
        pixel_data[174][71] = 1;
        pixel_data[174][72] = 1;
        pixel_data[174][73] = 1;
        pixel_data[174][74] = 1;
        pixel_data[174][75] = 1;
        pixel_data[174][76] = 1;
        pixel_data[174][77] = 1;
        pixel_data[174][78] = 1;
        pixel_data[174][79] = 1;
        pixel_data[174][80] = 1;
        pixel_data[174][81] = 1;
        pixel_data[174][82] = 1;
        pixel_data[174][83] = 1;
        pixel_data[174][84] = 1;
        pixel_data[174][85] = 1;
        pixel_data[174][86] = 1;
        pixel_data[174][87] = 1;
        pixel_data[174][88] = 1;
        pixel_data[174][89] = 1;
        pixel_data[174][90] = 1;
        pixel_data[174][91] = 1;
        pixel_data[174][92] = 1;
        pixel_data[174][93] = 1;
        pixel_data[174][94] = 1;
        pixel_data[174][95] = 1;
        pixel_data[174][96] = 1;
        pixel_data[174][97] = 1;
        pixel_data[174][98] = 1;
        pixel_data[174][99] = 1;
        pixel_data[174][100] = 1;
        pixel_data[174][101] = 1;
        pixel_data[174][102] = 1;
        pixel_data[174][103] = 1;
        pixel_data[174][104] = 1;
        pixel_data[174][105] = 1;
        pixel_data[174][106] = 1;
        pixel_data[174][107] = 1;
        pixel_data[174][108] = 1;
        pixel_data[174][109] = 1;
        pixel_data[174][110] = 1;
        pixel_data[174][111] = 1;
        pixel_data[174][112] = 1;
        pixel_data[174][113] = 1;
        pixel_data[174][114] = 1;
        pixel_data[174][115] = 1;
        pixel_data[174][116] = 1;
        pixel_data[174][117] = 1;
        pixel_data[174][118] = 5;
        pixel_data[174][119] = 7;
        pixel_data[174][120] = 10;
        pixel_data[174][121] = 12;
        pixel_data[174][122] = 13;
        pixel_data[174][123] = 13;
        pixel_data[174][124] = 13;
        pixel_data[174][125] = 13;
        pixel_data[174][126] = 13;
        pixel_data[174][127] = 13;
        pixel_data[174][128] = 13;
        pixel_data[174][129] = 10;
        pixel_data[174][130] = 7;
        pixel_data[174][131] = 2;
        pixel_data[174][132] = 1;
        pixel_data[174][133] = 1;
        pixel_data[174][134] = 1;
        pixel_data[174][135] = 1;
        pixel_data[174][136] = 1;
        pixel_data[174][137] = 1;
        pixel_data[174][138] = 1;
        pixel_data[174][139] = 1;
        pixel_data[174][140] = 1;
        pixel_data[174][141] = 1;
        pixel_data[174][142] = 1;
        pixel_data[174][143] = 1;
        pixel_data[174][144] = 1;
        pixel_data[174][145] = 1;
        pixel_data[174][146] = 1;
        pixel_data[174][147] = 1;
        pixel_data[174][148] = 1;
        pixel_data[174][149] = 1;
        pixel_data[174][150] = 1;
        pixel_data[174][151] = 1;
        pixel_data[174][152] = 1;
        pixel_data[174][153] = 1;
        pixel_data[174][154] = 1;
        pixel_data[174][155] = 1;
        pixel_data[174][156] = 1;
        pixel_data[174][157] = 1;
        pixel_data[174][158] = 1;
        pixel_data[174][159] = 1;
        pixel_data[174][160] = 1;
        pixel_data[174][161] = 1;
        pixel_data[174][162] = 1;
        pixel_data[174][163] = 1;
        pixel_data[174][164] = 1;
        pixel_data[174][165] = 1;
        pixel_data[174][166] = 1;
        pixel_data[174][167] = 1;
        pixel_data[174][168] = 1;
        pixel_data[174][169] = 1;
        pixel_data[174][170] = 1;
        pixel_data[174][171] = 1;
        pixel_data[174][172] = 1;
        pixel_data[174][173] = 1;
        pixel_data[174][174] = 1;
        pixel_data[174][175] = 1;
        pixel_data[174][176] = 1;
        pixel_data[174][177] = 1;
        pixel_data[174][178] = 1;
        pixel_data[174][179] = 1;
        pixel_data[174][180] = 1;
        pixel_data[174][181] = 1;
        pixel_data[174][182] = 1;
        pixel_data[174][183] = 1;
        pixel_data[174][184] = 6;
        pixel_data[174][185] = 9;
        pixel_data[174][186] = 11;
        pixel_data[174][187] = 11;
        pixel_data[174][188] = 0;
        pixel_data[174][189] = 0;
        pixel_data[174][190] = 0;
        pixel_data[174][191] = 0;
        pixel_data[174][192] = 0;
        pixel_data[174][193] = 0;
        pixel_data[174][194] = 0;
        pixel_data[174][195] = 0;
        pixel_data[174][196] = 0;
        pixel_data[174][197] = 0;
        pixel_data[174][198] = 0;
        pixel_data[174][199] = 0; // y=174
        pixel_data[175][0] = 0;
        pixel_data[175][1] = 0;
        pixel_data[175][2] = 0;
        pixel_data[175][3] = 0;
        pixel_data[175][4] = 0;
        pixel_data[175][5] = 11;
        pixel_data[175][6] = 11;
        pixel_data[175][7] = 8;
        pixel_data[175][8] = 4;
        pixel_data[175][9] = 1;
        pixel_data[175][10] = 1;
        pixel_data[175][11] = 1;
        pixel_data[175][12] = 4;
        pixel_data[175][13] = 4;
        pixel_data[175][14] = 2;
        pixel_data[175][15] = 1;
        pixel_data[175][16] = 1;
        pixel_data[175][17] = 1;
        pixel_data[175][18] = 1;
        pixel_data[175][19] = 1;
        pixel_data[175][20] = 1;
        pixel_data[175][21] = 1;
        pixel_data[175][22] = 1;
        pixel_data[175][23] = 1;
        pixel_data[175][24] = 1;
        pixel_data[175][25] = 1;
        pixel_data[175][26] = 1;
        pixel_data[175][27] = 1;
        pixel_data[175][28] = 1;
        pixel_data[175][29] = 1;
        pixel_data[175][30] = 1;
        pixel_data[175][31] = 1;
        pixel_data[175][32] = 1;
        pixel_data[175][33] = 1;
        pixel_data[175][34] = 1;
        pixel_data[175][35] = 1;
        pixel_data[175][36] = 1;
        pixel_data[175][37] = 1;
        pixel_data[175][38] = 1;
        pixel_data[175][39] = 1;
        pixel_data[175][40] = 1;
        pixel_data[175][41] = 1;
        pixel_data[175][42] = 1;
        pixel_data[175][43] = 1;
        pixel_data[175][44] = 1;
        pixel_data[175][45] = 1;
        pixel_data[175][46] = 1;
        pixel_data[175][47] = 1;
        pixel_data[175][48] = 1;
        pixel_data[175][49] = 1;
        pixel_data[175][50] = 1;
        pixel_data[175][51] = 1;
        pixel_data[175][52] = 1;
        pixel_data[175][53] = 1;
        pixel_data[175][54] = 1;
        pixel_data[175][55] = 1;
        pixel_data[175][56] = 1;
        pixel_data[175][57] = 1;
        pixel_data[175][58] = 1;
        pixel_data[175][59] = 1;
        pixel_data[175][60] = 1;
        pixel_data[175][61] = 1;
        pixel_data[175][62] = 1;
        pixel_data[175][63] = 1;
        pixel_data[175][64] = 1;
        pixel_data[175][65] = 1;
        pixel_data[175][66] = 1;
        pixel_data[175][67] = 1;
        pixel_data[175][68] = 1;
        pixel_data[175][69] = 1;
        pixel_data[175][70] = 1;
        pixel_data[175][71] = 1;
        pixel_data[175][72] = 1;
        pixel_data[175][73] = 1;
        pixel_data[175][74] = 1;
        pixel_data[175][75] = 1;
        pixel_data[175][76] = 1;
        pixel_data[175][77] = 1;
        pixel_data[175][78] = 1;
        pixel_data[175][79] = 1;
        pixel_data[175][80] = 1;
        pixel_data[175][81] = 1;
        pixel_data[175][82] = 1;
        pixel_data[175][83] = 1;
        pixel_data[175][84] = 1;
        pixel_data[175][85] = 1;
        pixel_data[175][86] = 1;
        pixel_data[175][87] = 1;
        pixel_data[175][88] = 1;
        pixel_data[175][89] = 1;
        pixel_data[175][90] = 1;
        pixel_data[175][91] = 1;
        pixel_data[175][92] = 1;
        pixel_data[175][93] = 1;
        pixel_data[175][94] = 1;
        pixel_data[175][95] = 1;
        pixel_data[175][96] = 1;
        pixel_data[175][97] = 1;
        pixel_data[175][98] = 1;
        pixel_data[175][99] = 1;
        pixel_data[175][100] = 1;
        pixel_data[175][101] = 1;
        pixel_data[175][102] = 1;
        pixel_data[175][103] = 1;
        pixel_data[175][104] = 1;
        pixel_data[175][105] = 1;
        pixel_data[175][106] = 1;
        pixel_data[175][107] = 1;
        pixel_data[175][108] = 1;
        pixel_data[175][109] = 1;
        pixel_data[175][110] = 1;
        pixel_data[175][111] = 1;
        pixel_data[175][112] = 1;
        pixel_data[175][113] = 1;
        pixel_data[175][114] = 1;
        pixel_data[175][115] = 4;
        pixel_data[175][116] = 8;
        pixel_data[175][117] = 12;
        pixel_data[175][118] = 13;
        pixel_data[175][119] = 13;
        pixel_data[175][120] = 13;
        pixel_data[175][121] = 13;
        pixel_data[175][122] = 13;
        pixel_data[175][123] = 13;
        pixel_data[175][124] = 13;
        pixel_data[175][125] = 13;
        pixel_data[175][126] = 13;
        pixel_data[175][127] = 13;
        pixel_data[175][128] = 13;
        pixel_data[175][129] = 13;
        pixel_data[175][130] = 13;
        pixel_data[175][131] = 13;
        pixel_data[175][132] = 12;
        pixel_data[175][133] = 6;
        pixel_data[175][134] = 1;
        pixel_data[175][135] = 1;
        pixel_data[175][136] = 1;
        pixel_data[175][137] = 1;
        pixel_data[175][138] = 1;
        pixel_data[175][139] = 1;
        pixel_data[175][140] = 1;
        pixel_data[175][141] = 1;
        pixel_data[175][142] = 1;
        pixel_data[175][143] = 1;
        pixel_data[175][144] = 1;
        pixel_data[175][145] = 1;
        pixel_data[175][146] = 1;
        pixel_data[175][147] = 1;
        pixel_data[175][148] = 1;
        pixel_data[175][149] = 1;
        pixel_data[175][150] = 1;
        pixel_data[175][151] = 1;
        pixel_data[175][152] = 1;
        pixel_data[175][153] = 1;
        pixel_data[175][154] = 1;
        pixel_data[175][155] = 1;
        pixel_data[175][156] = 1;
        pixel_data[175][157] = 1;
        pixel_data[175][158] = 1;
        pixel_data[175][159] = 1;
        pixel_data[175][160] = 1;
        pixel_data[175][161] = 1;
        pixel_data[175][162] = 1;
        pixel_data[175][163] = 1;
        pixel_data[175][164] = 1;
        pixel_data[175][165] = 1;
        pixel_data[175][166] = 1;
        pixel_data[175][167] = 1;
        pixel_data[175][168] = 1;
        pixel_data[175][169] = 1;
        pixel_data[175][170] = 1;
        pixel_data[175][171] = 1;
        pixel_data[175][172] = 1;
        pixel_data[175][173] = 1;
        pixel_data[175][174] = 1;
        pixel_data[175][175] = 1;
        pixel_data[175][176] = 1;
        pixel_data[175][177] = 1;
        pixel_data[175][178] = 1;
        pixel_data[175][179] = 1;
        pixel_data[175][180] = 1;
        pixel_data[175][181] = 1;
        pixel_data[175][182] = 1;
        pixel_data[175][183] = 1;
        pixel_data[175][184] = 1;
        pixel_data[175][185] = 6;
        pixel_data[175][186] = 9;
        pixel_data[175][187] = 11;
        pixel_data[175][188] = 11;
        pixel_data[175][189] = 0;
        pixel_data[175][190] = 0;
        pixel_data[175][191] = 0;
        pixel_data[175][192] = 0;
        pixel_data[175][193] = 0;
        pixel_data[175][194] = 0;
        pixel_data[175][195] = 0;
        pixel_data[175][196] = 0;
        pixel_data[175][197] = 0;
        pixel_data[175][198] = 0;
        pixel_data[175][199] = 0; // y=175
        pixel_data[176][0] = 0;
        pixel_data[176][1] = 0;
        pixel_data[176][2] = 0;
        pixel_data[176][3] = 0;
        pixel_data[176][4] = 0;
        pixel_data[176][5] = 11;
        pixel_data[176][6] = 11;
        pixel_data[176][7] = 8;
        pixel_data[176][8] = 4;
        pixel_data[176][9] = 1;
        pixel_data[176][10] = 1;
        pixel_data[176][11] = 1;
        pixel_data[176][12] = 4;
        pixel_data[176][13] = 4;
        pixel_data[176][14] = 2;
        pixel_data[176][15] = 1;
        pixel_data[176][16] = 1;
        pixel_data[176][17] = 1;
        pixel_data[176][18] = 1;
        pixel_data[176][19] = 1;
        pixel_data[176][20] = 1;
        pixel_data[176][21] = 1;
        pixel_data[176][22] = 1;
        pixel_data[176][23] = 1;
        pixel_data[176][24] = 1;
        pixel_data[176][25] = 1;
        pixel_data[176][26] = 1;
        pixel_data[176][27] = 1;
        pixel_data[176][28] = 1;
        pixel_data[176][29] = 1;
        pixel_data[176][30] = 1;
        pixel_data[176][31] = 1;
        pixel_data[176][32] = 1;
        pixel_data[176][33] = 1;
        pixel_data[176][34] = 1;
        pixel_data[176][35] = 1;
        pixel_data[176][36] = 1;
        pixel_data[176][37] = 1;
        pixel_data[176][38] = 1;
        pixel_data[176][39] = 1;
        pixel_data[176][40] = 1;
        pixel_data[176][41] = 1;
        pixel_data[176][42] = 1;
        pixel_data[176][43] = 1;
        pixel_data[176][44] = 1;
        pixel_data[176][45] = 1;
        pixel_data[176][46] = 1;
        pixel_data[176][47] = 1;
        pixel_data[176][48] = 1;
        pixel_data[176][49] = 1;
        pixel_data[176][50] = 1;
        pixel_data[176][51] = 1;
        pixel_data[176][52] = 1;
        pixel_data[176][53] = 1;
        pixel_data[176][54] = 1;
        pixel_data[176][55] = 1;
        pixel_data[176][56] = 1;
        pixel_data[176][57] = 1;
        pixel_data[176][58] = 1;
        pixel_data[176][59] = 1;
        pixel_data[176][60] = 1;
        pixel_data[176][61] = 1;
        pixel_data[176][62] = 1;
        pixel_data[176][63] = 1;
        pixel_data[176][64] = 1;
        pixel_data[176][65] = 1;
        pixel_data[176][66] = 1;
        pixel_data[176][67] = 1;
        pixel_data[176][68] = 1;
        pixel_data[176][69] = 1;
        pixel_data[176][70] = 1;
        pixel_data[176][71] = 1;
        pixel_data[176][72] = 1;
        pixel_data[176][73] = 1;
        pixel_data[176][74] = 1;
        pixel_data[176][75] = 1;
        pixel_data[176][76] = 1;
        pixel_data[176][77] = 1;
        pixel_data[176][78] = 1;
        pixel_data[176][79] = 1;
        pixel_data[176][80] = 1;
        pixel_data[176][81] = 1;
        pixel_data[176][82] = 1;
        pixel_data[176][83] = 1;
        pixel_data[176][84] = 1;
        pixel_data[176][85] = 1;
        pixel_data[176][86] = 1;
        pixel_data[176][87] = 1;
        pixel_data[176][88] = 1;
        pixel_data[176][89] = 1;
        pixel_data[176][90] = 1;
        pixel_data[176][91] = 1;
        pixel_data[176][92] = 1;
        pixel_data[176][93] = 1;
        pixel_data[176][94] = 1;
        pixel_data[176][95] = 1;
        pixel_data[176][96] = 1;
        pixel_data[176][97] = 1;
        pixel_data[176][98] = 1;
        pixel_data[176][99] = 1;
        pixel_data[176][100] = 1;
        pixel_data[176][101] = 1;
        pixel_data[176][102] = 1;
        pixel_data[176][103] = 1;
        pixel_data[176][104] = 1;
        pixel_data[176][105] = 1;
        pixel_data[176][106] = 1;
        pixel_data[176][107] = 1;
        pixel_data[176][108] = 1;
        pixel_data[176][109] = 1;
        pixel_data[176][110] = 1;
        pixel_data[176][111] = 1;
        pixel_data[176][112] = 1;
        pixel_data[176][113] = 1;
        pixel_data[176][114] = 6;
        pixel_data[176][115] = 10;
        pixel_data[176][116] = 13;
        pixel_data[176][117] = 13;
        pixel_data[176][118] = 13;
        pixel_data[176][119] = 13;
        pixel_data[176][120] = 13;
        pixel_data[176][121] = 13;
        pixel_data[176][122] = 13;
        pixel_data[176][123] = 13;
        pixel_data[176][124] = 13;
        pixel_data[176][125] = 13;
        pixel_data[176][126] = 13;
        pixel_data[176][127] = 13;
        pixel_data[176][128] = 13;
        pixel_data[176][129] = 13;
        pixel_data[176][130] = 13;
        pixel_data[176][131] = 13;
        pixel_data[176][132] = 13;
        pixel_data[176][133] = 13;
        pixel_data[176][134] = 9;
        pixel_data[176][135] = 4;
        pixel_data[176][136] = 1;
        pixel_data[176][137] = 1;
        pixel_data[176][138] = 1;
        pixel_data[176][139] = 1;
        pixel_data[176][140] = 1;
        pixel_data[176][141] = 1;
        pixel_data[176][142] = 1;
        pixel_data[176][143] = 1;
        pixel_data[176][144] = 1;
        pixel_data[176][145] = 1;
        pixel_data[176][146] = 1;
        pixel_data[176][147] = 1;
        pixel_data[176][148] = 1;
        pixel_data[176][149] = 1;
        pixel_data[176][150] = 1;
        pixel_data[176][151] = 1;
        pixel_data[176][152] = 1;
        pixel_data[176][153] = 1;
        pixel_data[176][154] = 1;
        pixel_data[176][155] = 1;
        pixel_data[176][156] = 1;
        pixel_data[176][157] = 1;
        pixel_data[176][158] = 1;
        pixel_data[176][159] = 1;
        pixel_data[176][160] = 1;
        pixel_data[176][161] = 1;
        pixel_data[176][162] = 1;
        pixel_data[176][163] = 1;
        pixel_data[176][164] = 1;
        pixel_data[176][165] = 1;
        pixel_data[176][166] = 1;
        pixel_data[176][167] = 1;
        pixel_data[176][168] = 1;
        pixel_data[176][169] = 1;
        pixel_data[176][170] = 1;
        pixel_data[176][171] = 1;
        pixel_data[176][172] = 1;
        pixel_data[176][173] = 1;
        pixel_data[176][174] = 1;
        pixel_data[176][175] = 1;
        pixel_data[176][176] = 1;
        pixel_data[176][177] = 1;
        pixel_data[176][178] = 1;
        pixel_data[176][179] = 1;
        pixel_data[176][180] = 1;
        pixel_data[176][181] = 1;
        pixel_data[176][182] = 1;
        pixel_data[176][183] = 1;
        pixel_data[176][184] = 1;
        pixel_data[176][185] = 4;
        pixel_data[176][186] = 7;
        pixel_data[176][187] = 9;
        pixel_data[176][188] = 11;
        pixel_data[176][189] = 13;
        pixel_data[176][190] = 0;
        pixel_data[176][191] = 0;
        pixel_data[176][192] = 0;
        pixel_data[176][193] = 0;
        pixel_data[176][194] = 0;
        pixel_data[176][195] = 0;
        pixel_data[176][196] = 0;
        pixel_data[176][197] = 0;
        pixel_data[176][198] = 0;
        pixel_data[176][199] = 0; // y=176
        pixel_data[177][0] = 0;
        pixel_data[177][1] = 0;
        pixel_data[177][2] = 0;
        pixel_data[177][3] = 0;
        pixel_data[177][4] = 11;
        pixel_data[177][5] = 11;
        pixel_data[177][6] = 11;
        pixel_data[177][7] = 7;
        pixel_data[177][8] = 1;
        pixel_data[177][9] = 1;
        pixel_data[177][10] = 1;
        pixel_data[177][11] = 1;
        pixel_data[177][12] = 4;
        pixel_data[177][13] = 4;
        pixel_data[177][14] = 2;
        pixel_data[177][15] = 1;
        pixel_data[177][16] = 1;
        pixel_data[177][17] = 1;
        pixel_data[177][18] = 1;
        pixel_data[177][19] = 1;
        pixel_data[177][20] = 1;
        pixel_data[177][21] = 1;
        pixel_data[177][22] = 1;
        pixel_data[177][23] = 1;
        pixel_data[177][24] = 1;
        pixel_data[177][25] = 1;
        pixel_data[177][26] = 1;
        pixel_data[177][27] = 1;
        pixel_data[177][28] = 1;
        pixel_data[177][29] = 1;
        pixel_data[177][30] = 1;
        pixel_data[177][31] = 1;
        pixel_data[177][32] = 1;
        pixel_data[177][33] = 1;
        pixel_data[177][34] = 1;
        pixel_data[177][35] = 1;
        pixel_data[177][36] = 1;
        pixel_data[177][37] = 1;
        pixel_data[177][38] = 1;
        pixel_data[177][39] = 1;
        pixel_data[177][40] = 1;
        pixel_data[177][41] = 1;
        pixel_data[177][42] = 1;
        pixel_data[177][43] = 1;
        pixel_data[177][44] = 1;
        pixel_data[177][45] = 1;
        pixel_data[177][46] = 1;
        pixel_data[177][47] = 1;
        pixel_data[177][48] = 1;
        pixel_data[177][49] = 1;
        pixel_data[177][50] = 1;
        pixel_data[177][51] = 1;
        pixel_data[177][52] = 1;
        pixel_data[177][53] = 1;
        pixel_data[177][54] = 1;
        pixel_data[177][55] = 1;
        pixel_data[177][56] = 1;
        pixel_data[177][57] = 1;
        pixel_data[177][58] = 1;
        pixel_data[177][59] = 1;
        pixel_data[177][60] = 1;
        pixel_data[177][61] = 1;
        pixel_data[177][62] = 1;
        pixel_data[177][63] = 1;
        pixel_data[177][64] = 1;
        pixel_data[177][65] = 1;
        pixel_data[177][66] = 1;
        pixel_data[177][67] = 1;
        pixel_data[177][68] = 1;
        pixel_data[177][69] = 1;
        pixel_data[177][70] = 1;
        pixel_data[177][71] = 1;
        pixel_data[177][72] = 1;
        pixel_data[177][73] = 1;
        pixel_data[177][74] = 1;
        pixel_data[177][75] = 1;
        pixel_data[177][76] = 1;
        pixel_data[177][77] = 1;
        pixel_data[177][78] = 1;
        pixel_data[177][79] = 1;
        pixel_data[177][80] = 1;
        pixel_data[177][81] = 1;
        pixel_data[177][82] = 1;
        pixel_data[177][83] = 1;
        pixel_data[177][84] = 1;
        pixel_data[177][85] = 1;
        pixel_data[177][86] = 1;
        pixel_data[177][87] = 1;
        pixel_data[177][88] = 1;
        pixel_data[177][89] = 1;
        pixel_data[177][90] = 1;
        pixel_data[177][91] = 1;
        pixel_data[177][92] = 1;
        pixel_data[177][93] = 1;
        pixel_data[177][94] = 1;
        pixel_data[177][95] = 1;
        pixel_data[177][96] = 1;
        pixel_data[177][97] = 1;
        pixel_data[177][98] = 1;
        pixel_data[177][99] = 1;
        pixel_data[177][100] = 1;
        pixel_data[177][101] = 1;
        pixel_data[177][102] = 1;
        pixel_data[177][103] = 1;
        pixel_data[177][104] = 1;
        pixel_data[177][105] = 1;
        pixel_data[177][106] = 1;
        pixel_data[177][107] = 1;
        pixel_data[177][108] = 1;
        pixel_data[177][109] = 1;
        pixel_data[177][110] = 1;
        pixel_data[177][111] = 1;
        pixel_data[177][112] = 1;
        pixel_data[177][113] = 6;
        pixel_data[177][114] = 10;
        pixel_data[177][115] = 13;
        pixel_data[177][116] = 13;
        pixel_data[177][117] = 13;
        pixel_data[177][118] = 13;
        pixel_data[177][119] = 13;
        pixel_data[177][120] = 13;
        pixel_data[177][121] = 13;
        pixel_data[177][122] = 13;
        pixel_data[177][123] = 13;
        pixel_data[177][124] = 13;
        pixel_data[177][125] = 13;
        pixel_data[177][126] = 13;
        pixel_data[177][127] = 13;
        pixel_data[177][128] = 13;
        pixel_data[177][129] = 13;
        pixel_data[177][130] = 13;
        pixel_data[177][131] = 13;
        pixel_data[177][132] = 13;
        pixel_data[177][133] = 13;
        pixel_data[177][134] = 13;
        pixel_data[177][135] = 10;
        pixel_data[177][136] = 5;
        pixel_data[177][137] = 1;
        pixel_data[177][138] = 1;
        pixel_data[177][139] = 1;
        pixel_data[177][140] = 1;
        pixel_data[177][141] = 1;
        pixel_data[177][142] = 1;
        pixel_data[177][143] = 1;
        pixel_data[177][144] = 1;
        pixel_data[177][145] = 1;
        pixel_data[177][146] = 1;
        pixel_data[177][147] = 1;
        pixel_data[177][148] = 1;
        pixel_data[177][149] = 1;
        pixel_data[177][150] = 1;
        pixel_data[177][151] = 1;
        pixel_data[177][152] = 1;
        pixel_data[177][153] = 1;
        pixel_data[177][154] = 1;
        pixel_data[177][155] = 1;
        pixel_data[177][156] = 1;
        pixel_data[177][157] = 1;
        pixel_data[177][158] = 1;
        pixel_data[177][159] = 1;
        pixel_data[177][160] = 1;
        pixel_data[177][161] = 1;
        pixel_data[177][162] = 1;
        pixel_data[177][163] = 1;
        pixel_data[177][164] = 1;
        pixel_data[177][165] = 1;
        pixel_data[177][166] = 1;
        pixel_data[177][167] = 1;
        pixel_data[177][168] = 1;
        pixel_data[177][169] = 1;
        pixel_data[177][170] = 1;
        pixel_data[177][171] = 1;
        pixel_data[177][172] = 1;
        pixel_data[177][173] = 1;
        pixel_data[177][174] = 1;
        pixel_data[177][175] = 1;
        pixel_data[177][176] = 1;
        pixel_data[177][177] = 1;
        pixel_data[177][178] = 1;
        pixel_data[177][179] = 1;
        pixel_data[177][180] = 1;
        pixel_data[177][181] = 1;
        pixel_data[177][182] = 1;
        pixel_data[177][183] = 1;
        pixel_data[177][184] = 1;
        pixel_data[177][185] = 1;
        pixel_data[177][186] = 6;
        pixel_data[177][187] = 8;
        pixel_data[177][188] = 11;
        pixel_data[177][189] = 11;
        pixel_data[177][190] = 0;
        pixel_data[177][191] = 0;
        pixel_data[177][192] = 0;
        pixel_data[177][193] = 0;
        pixel_data[177][194] = 0;
        pixel_data[177][195] = 0;
        pixel_data[177][196] = 0;
        pixel_data[177][197] = 0;
        pixel_data[177][198] = 0;
        pixel_data[177][199] = 0; // y=177
        pixel_data[178][0] = 0;
        pixel_data[178][1] = 0;
        pixel_data[178][2] = 0;
        pixel_data[178][3] = 0;
        pixel_data[178][4] = 11;
        pixel_data[178][5] = 11;
        pixel_data[178][6] = 11;
        pixel_data[178][7] = 7;
        pixel_data[178][8] = 1;
        pixel_data[178][9] = 1;
        pixel_data[178][10] = 1;
        pixel_data[178][11] = 1;
        pixel_data[178][12] = 4;
        pixel_data[178][13] = 4;
        pixel_data[178][14] = 2;
        pixel_data[178][15] = 1;
        pixel_data[178][16] = 1;
        pixel_data[178][17] = 1;
        pixel_data[178][18] = 1;
        pixel_data[178][19] = 1;
        pixel_data[178][20] = 1;
        pixel_data[178][21] = 1;
        pixel_data[178][22] = 1;
        pixel_data[178][23] = 1;
        pixel_data[178][24] = 1;
        pixel_data[178][25] = 1;
        pixel_data[178][26] = 1;
        pixel_data[178][27] = 1;
        pixel_data[178][28] = 1;
        pixel_data[178][29] = 1;
        pixel_data[178][30] = 1;
        pixel_data[178][31] = 1;
        pixel_data[178][32] = 1;
        pixel_data[178][33] = 1;
        pixel_data[178][34] = 1;
        pixel_data[178][35] = 1;
        pixel_data[178][36] = 1;
        pixel_data[178][37] = 1;
        pixel_data[178][38] = 1;
        pixel_data[178][39] = 1;
        pixel_data[178][40] = 1;
        pixel_data[178][41] = 1;
        pixel_data[178][42] = 1;
        pixel_data[178][43] = 1;
        pixel_data[178][44] = 1;
        pixel_data[178][45] = 1;
        pixel_data[178][46] = 1;
        pixel_data[178][47] = 1;
        pixel_data[178][48] = 1;
        pixel_data[178][49] = 1;
        pixel_data[178][50] = 1;
        pixel_data[178][51] = 1;
        pixel_data[178][52] = 1;
        pixel_data[178][53] = 1;
        pixel_data[178][54] = 1;
        pixel_data[178][55] = 1;
        pixel_data[178][56] = 1;
        pixel_data[178][57] = 1;
        pixel_data[178][58] = 1;
        pixel_data[178][59] = 1;
        pixel_data[178][60] = 1;
        pixel_data[178][61] = 1;
        pixel_data[178][62] = 1;
        pixel_data[178][63] = 1;
        pixel_data[178][64] = 1;
        pixel_data[178][65] = 1;
        pixel_data[178][66] = 1;
        pixel_data[178][67] = 1;
        pixel_data[178][68] = 1;
        pixel_data[178][69] = 1;
        pixel_data[178][70] = 1;
        pixel_data[178][71] = 1;
        pixel_data[178][72] = 1;
        pixel_data[178][73] = 1;
        pixel_data[178][74] = 1;
        pixel_data[178][75] = 1;
        pixel_data[178][76] = 1;
        pixel_data[178][77] = 1;
        pixel_data[178][78] = 1;
        pixel_data[178][79] = 1;
        pixel_data[178][80] = 1;
        pixel_data[178][81] = 1;
        pixel_data[178][82] = 1;
        pixel_data[178][83] = 1;
        pixel_data[178][84] = 1;
        pixel_data[178][85] = 1;
        pixel_data[178][86] = 1;
        pixel_data[178][87] = 1;
        pixel_data[178][88] = 1;
        pixel_data[178][89] = 1;
        pixel_data[178][90] = 1;
        pixel_data[178][91] = 1;
        pixel_data[178][92] = 1;
        pixel_data[178][93] = 1;
        pixel_data[178][94] = 1;
        pixel_data[178][95] = 1;
        pixel_data[178][96] = 1;
        pixel_data[178][97] = 1;
        pixel_data[178][98] = 1;
        pixel_data[178][99] = 1;
        pixel_data[178][100] = 1;
        pixel_data[178][101] = 1;
        pixel_data[178][102] = 1;
        pixel_data[178][103] = 1;
        pixel_data[178][104] = 1;
        pixel_data[178][105] = 1;
        pixel_data[178][106] = 1;
        pixel_data[178][107] = 1;
        pixel_data[178][108] = 1;
        pixel_data[178][109] = 1;
        pixel_data[178][110] = 1;
        pixel_data[178][111] = 1;
        pixel_data[178][112] = 5;
        pixel_data[178][113] = 9;
        pixel_data[178][114] = 13;
        pixel_data[178][115] = 13;
        pixel_data[178][116] = 13;
        pixel_data[178][117] = 13;
        pixel_data[178][118] = 13;
        pixel_data[178][119] = 13;
        pixel_data[178][120] = 13;
        pixel_data[178][121] = 13;
        pixel_data[178][122] = 13;
        pixel_data[178][123] = 13;
        pixel_data[178][124] = 13;
        pixel_data[178][125] = 13;
        pixel_data[178][126] = 13;
        pixel_data[178][127] = 13;
        pixel_data[178][128] = 13;
        pixel_data[178][129] = 13;
        pixel_data[178][130] = 13;
        pixel_data[178][131] = 13;
        pixel_data[178][132] = 13;
        pixel_data[178][133] = 13;
        pixel_data[178][134] = 13;
        pixel_data[178][135] = 13;
        pixel_data[178][136] = 9;
        pixel_data[178][137] = 4;
        pixel_data[178][138] = 1;
        pixel_data[178][139] = 1;
        pixel_data[178][140] = 1;
        pixel_data[178][141] = 1;
        pixel_data[178][142] = 1;
        pixel_data[178][143] = 1;
        pixel_data[178][144] = 1;
        pixel_data[178][145] = 1;
        pixel_data[178][146] = 1;
        pixel_data[178][147] = 1;
        pixel_data[178][148] = 1;
        pixel_data[178][149] = 1;
        pixel_data[178][150] = 1;
        pixel_data[178][151] = 1;
        pixel_data[178][152] = 1;
        pixel_data[178][153] = 1;
        pixel_data[178][154] = 1;
        pixel_data[178][155] = 1;
        pixel_data[178][156] = 1;
        pixel_data[178][157] = 1;
        pixel_data[178][158] = 1;
        pixel_data[178][159] = 1;
        pixel_data[178][160] = 1;
        pixel_data[178][161] = 1;
        pixel_data[178][162] = 1;
        pixel_data[178][163] = 1;
        pixel_data[178][164] = 1;
        pixel_data[178][165] = 1;
        pixel_data[178][166] = 1;
        pixel_data[178][167] = 1;
        pixel_data[178][168] = 1;
        pixel_data[178][169] = 1;
        pixel_data[178][170] = 1;
        pixel_data[178][171] = 1;
        pixel_data[178][172] = 1;
        pixel_data[178][173] = 1;
        pixel_data[178][174] = 1;
        pixel_data[178][175] = 1;
        pixel_data[178][176] = 1;
        pixel_data[178][177] = 1;
        pixel_data[178][178] = 1;
        pixel_data[178][179] = 1;
        pixel_data[178][180] = 1;
        pixel_data[178][181] = 1;
        pixel_data[178][182] = 1;
        pixel_data[178][183] = 1;
        pixel_data[178][184] = 1;
        pixel_data[178][185] = 1;
        pixel_data[178][186] = 4;
        pixel_data[178][187] = 7;
        pixel_data[178][188] = 11;
        pixel_data[178][189] = 11;
        pixel_data[178][190] = 0;
        pixel_data[178][191] = 0;
        pixel_data[178][192] = 0;
        pixel_data[178][193] = 0;
        pixel_data[178][194] = 0;
        pixel_data[178][195] = 0;
        pixel_data[178][196] = 0;
        pixel_data[178][197] = 0;
        pixel_data[178][198] = 0;
        pixel_data[178][199] = 0; // y=178
        pixel_data[179][0] = 0;
        pixel_data[179][1] = 0;
        pixel_data[179][2] = 0;
        pixel_data[179][3] = 0;
        pixel_data[179][4] = 11;
        pixel_data[179][5] = 11;
        pixel_data[179][6] = 11;
        pixel_data[179][7] = 7;
        pixel_data[179][8] = 1;
        pixel_data[179][9] = 1;
        pixel_data[179][10] = 1;
        pixel_data[179][11] = 1;
        pixel_data[179][12] = 4;
        pixel_data[179][13] = 4;
        pixel_data[179][14] = 2;
        pixel_data[179][15] = 1;
        pixel_data[179][16] = 1;
        pixel_data[179][17] = 1;
        pixel_data[179][18] = 1;
        pixel_data[179][19] = 1;
        pixel_data[179][20] = 1;
        pixel_data[179][21] = 1;
        pixel_data[179][22] = 1;
        pixel_data[179][23] = 1;
        pixel_data[179][24] = 1;
        pixel_data[179][25] = 1;
        pixel_data[179][26] = 1;
        pixel_data[179][27] = 1;
        pixel_data[179][28] = 1;
        pixel_data[179][29] = 1;
        pixel_data[179][30] = 1;
        pixel_data[179][31] = 1;
        pixel_data[179][32] = 1;
        pixel_data[179][33] = 1;
        pixel_data[179][34] = 1;
        pixel_data[179][35] = 1;
        pixel_data[179][36] = 1;
        pixel_data[179][37] = 1;
        pixel_data[179][38] = 1;
        pixel_data[179][39] = 1;
        pixel_data[179][40] = 1;
        pixel_data[179][41] = 1;
        pixel_data[179][42] = 1;
        pixel_data[179][43] = 1;
        pixel_data[179][44] = 1;
        pixel_data[179][45] = 1;
        pixel_data[179][46] = 1;
        pixel_data[179][47] = 1;
        pixel_data[179][48] = 1;
        pixel_data[179][49] = 1;
        pixel_data[179][50] = 1;
        pixel_data[179][51] = 1;
        pixel_data[179][52] = 1;
        pixel_data[179][53] = 1;
        pixel_data[179][54] = 1;
        pixel_data[179][55] = 1;
        pixel_data[179][56] = 1;
        pixel_data[179][57] = 1;
        pixel_data[179][58] = 1;
        pixel_data[179][59] = 1;
        pixel_data[179][60] = 1;
        pixel_data[179][61] = 1;
        pixel_data[179][62] = 1;
        pixel_data[179][63] = 1;
        pixel_data[179][64] = 1;
        pixel_data[179][65] = 1;
        pixel_data[179][66] = 1;
        pixel_data[179][67] = 1;
        pixel_data[179][68] = 1;
        pixel_data[179][69] = 1;
        pixel_data[179][70] = 1;
        pixel_data[179][71] = 1;
        pixel_data[179][72] = 1;
        pixel_data[179][73] = 1;
        pixel_data[179][74] = 1;
        pixel_data[179][75] = 1;
        pixel_data[179][76] = 1;
        pixel_data[179][77] = 1;
        pixel_data[179][78] = 1;
        pixel_data[179][79] = 1;
        pixel_data[179][80] = 1;
        pixel_data[179][81] = 1;
        pixel_data[179][82] = 1;
        pixel_data[179][83] = 1;
        pixel_data[179][84] = 1;
        pixel_data[179][85] = 1;
        pixel_data[179][86] = 1;
        pixel_data[179][87] = 1;
        pixel_data[179][88] = 1;
        pixel_data[179][89] = 1;
        pixel_data[179][90] = 1;
        pixel_data[179][91] = 1;
        pixel_data[179][92] = 1;
        pixel_data[179][93] = 1;
        pixel_data[179][94] = 1;
        pixel_data[179][95] = 1;
        pixel_data[179][96] = 1;
        pixel_data[179][97] = 1;
        pixel_data[179][98] = 1;
        pixel_data[179][99] = 1;
        pixel_data[179][100] = 1;
        pixel_data[179][101] = 1;
        pixel_data[179][102] = 1;
        pixel_data[179][103] = 1;
        pixel_data[179][104] = 1;
        pixel_data[179][105] = 1;
        pixel_data[179][106] = 1;
        pixel_data[179][107] = 1;
        pixel_data[179][108] = 1;
        pixel_data[179][109] = 1;
        pixel_data[179][110] = 1;
        pixel_data[179][111] = 1;
        pixel_data[179][112] = 5;
        pixel_data[179][113] = 10;
        pixel_data[179][114] = 13;
        pixel_data[179][115] = 13;
        pixel_data[179][116] = 13;
        pixel_data[179][117] = 13;
        pixel_data[179][118] = 13;
        pixel_data[179][119] = 13;
        pixel_data[179][120] = 13;
        pixel_data[179][121] = 13;
        pixel_data[179][122] = 13;
        pixel_data[179][123] = 13;
        pixel_data[179][124] = 13;
        pixel_data[179][125] = 13;
        pixel_data[179][126] = 13;
        pixel_data[179][127] = 13;
        pixel_data[179][128] = 13;
        pixel_data[179][129] = 13;
        pixel_data[179][130] = 13;
        pixel_data[179][131] = 13;
        pixel_data[179][132] = 13;
        pixel_data[179][133] = 13;
        pixel_data[179][134] = 13;
        pixel_data[179][135] = 13;
        pixel_data[179][136] = 10;
        pixel_data[179][137] = 5;
        pixel_data[179][138] = 1;
        pixel_data[179][139] = 1;
        pixel_data[179][140] = 1;
        pixel_data[179][141] = 1;
        pixel_data[179][142] = 1;
        pixel_data[179][143] = 1;
        pixel_data[179][144] = 1;
        pixel_data[179][145] = 1;
        pixel_data[179][146] = 1;
        pixel_data[179][147] = 1;
        pixel_data[179][148] = 1;
        pixel_data[179][149] = 1;
        pixel_data[179][150] = 1;
        pixel_data[179][151] = 1;
        pixel_data[179][152] = 1;
        pixel_data[179][153] = 1;
        pixel_data[179][154] = 1;
        pixel_data[179][155] = 1;
        pixel_data[179][156] = 1;
        pixel_data[179][157] = 1;
        pixel_data[179][158] = 1;
        pixel_data[179][159] = 1;
        pixel_data[179][160] = 1;
        pixel_data[179][161] = 1;
        pixel_data[179][162] = 1;
        pixel_data[179][163] = 1;
        pixel_data[179][164] = 1;
        pixel_data[179][165] = 1;
        pixel_data[179][166] = 1;
        pixel_data[179][167] = 1;
        pixel_data[179][168] = 1;
        pixel_data[179][169] = 1;
        pixel_data[179][170] = 1;
        pixel_data[179][171] = 1;
        pixel_data[179][172] = 1;
        pixel_data[179][173] = 1;
        pixel_data[179][174] = 1;
        pixel_data[179][175] = 1;
        pixel_data[179][176] = 1;
        pixel_data[179][177] = 1;
        pixel_data[179][178] = 1;
        pixel_data[179][179] = 1;
        pixel_data[179][180] = 1;
        pixel_data[179][181] = 1;
        pixel_data[179][182] = 1;
        pixel_data[179][183] = 1;
        pixel_data[179][184] = 1;
        pixel_data[179][185] = 1;
        pixel_data[179][186] = 1;
        pixel_data[179][187] = 7;
        pixel_data[179][188] = 9;
        pixel_data[179][189] = 11;
        pixel_data[179][190] = 10;
        pixel_data[179][191] = 0;
        pixel_data[179][192] = 0;
        pixel_data[179][193] = 0;
        pixel_data[179][194] = 0;
        pixel_data[179][195] = 0;
        pixel_data[179][196] = 0;
        pixel_data[179][197] = 0;
        pixel_data[179][198] = 0;
        pixel_data[179][199] = 0; // y=179
        pixel_data[180][0] = 0;
        pixel_data[180][1] = 0;
        pixel_data[180][2] = 0;
        pixel_data[180][3] = 0;
        pixel_data[180][4] = 11;
        pixel_data[180][5] = 11;
        pixel_data[180][6] = 11;
        pixel_data[180][7] = 7;
        pixel_data[180][8] = 1;
        pixel_data[180][9] = 1;
        pixel_data[180][10] = 1;
        pixel_data[180][11] = 1;
        pixel_data[180][12] = 4;
        pixel_data[180][13] = 4;
        pixel_data[180][14] = 4;
        pixel_data[180][15] = 1;
        pixel_data[180][16] = 1;
        pixel_data[180][17] = 1;
        pixel_data[180][18] = 1;
        pixel_data[180][19] = 1;
        pixel_data[180][20] = 1;
        pixel_data[180][21] = 1;
        pixel_data[180][22] = 1;
        pixel_data[180][23] = 1;
        pixel_data[180][24] = 1;
        pixel_data[180][25] = 1;
        pixel_data[180][26] = 1;
        pixel_data[180][27] = 1;
        pixel_data[180][28] = 1;
        pixel_data[180][29] = 1;
        pixel_data[180][30] = 1;
        pixel_data[180][31] = 1;
        pixel_data[180][32] = 1;
        pixel_data[180][33] = 1;
        pixel_data[180][34] = 1;
        pixel_data[180][35] = 1;
        pixel_data[180][36] = 1;
        pixel_data[180][37] = 1;
        pixel_data[180][38] = 1;
        pixel_data[180][39] = 1;
        pixel_data[180][40] = 1;
        pixel_data[180][41] = 1;
        pixel_data[180][42] = 1;
        pixel_data[180][43] = 1;
        pixel_data[180][44] = 1;
        pixel_data[180][45] = 1;
        pixel_data[180][46] = 1;
        pixel_data[180][47] = 1;
        pixel_data[180][48] = 1;
        pixel_data[180][49] = 1;
        pixel_data[180][50] = 1;
        pixel_data[180][51] = 1;
        pixel_data[180][52] = 1;
        pixel_data[180][53] = 1;
        pixel_data[180][54] = 1;
        pixel_data[180][55] = 1;
        pixel_data[180][56] = 1;
        pixel_data[180][57] = 1;
        pixel_data[180][58] = 1;
        pixel_data[180][59] = 1;
        pixel_data[180][60] = 1;
        pixel_data[180][61] = 1;
        pixel_data[180][62] = 1;
        pixel_data[180][63] = 1;
        pixel_data[180][64] = 1;
        pixel_data[180][65] = 1;
        pixel_data[180][66] = 1;
        pixel_data[180][67] = 1;
        pixel_data[180][68] = 1;
        pixel_data[180][69] = 1;
        pixel_data[180][70] = 1;
        pixel_data[180][71] = 1;
        pixel_data[180][72] = 1;
        pixel_data[180][73] = 1;
        pixel_data[180][74] = 1;
        pixel_data[180][75] = 1;
        pixel_data[180][76] = 1;
        pixel_data[180][77] = 1;
        pixel_data[180][78] = 1;
        pixel_data[180][79] = 1;
        pixel_data[180][80] = 1;
        pixel_data[180][81] = 1;
        pixel_data[180][82] = 1;
        pixel_data[180][83] = 1;
        pixel_data[180][84] = 1;
        pixel_data[180][85] = 1;
        pixel_data[180][86] = 1;
        pixel_data[180][87] = 1;
        pixel_data[180][88] = 1;
        pixel_data[180][89] = 1;
        pixel_data[180][90] = 1;
        pixel_data[180][91] = 1;
        pixel_data[180][92] = 1;
        pixel_data[180][93] = 1;
        pixel_data[180][94] = 1;
        pixel_data[180][95] = 1;
        pixel_data[180][96] = 1;
        pixel_data[180][97] = 1;
        pixel_data[180][98] = 1;
        pixel_data[180][99] = 1;
        pixel_data[180][100] = 1;
        pixel_data[180][101] = 1;
        pixel_data[180][102] = 1;
        pixel_data[180][103] = 1;
        pixel_data[180][104] = 1;
        pixel_data[180][105] = 1;
        pixel_data[180][106] = 1;
        pixel_data[180][107] = 1;
        pixel_data[180][108] = 1;
        pixel_data[180][109] = 1;
        pixel_data[180][110] = 1;
        pixel_data[180][111] = 1;
        pixel_data[180][112] = 4;
        pixel_data[180][113] = 9;
        pixel_data[180][114] = 13;
        pixel_data[180][115] = 13;
        pixel_data[180][116] = 13;
        pixel_data[180][117] = 13;
        pixel_data[180][118] = 13;
        pixel_data[180][119] = 13;
        pixel_data[180][120] = 13;
        pixel_data[180][121] = 13;
        pixel_data[180][122] = 13;
        pixel_data[180][123] = 13;
        pixel_data[180][124] = 13;
        pixel_data[180][125] = 13;
        pixel_data[180][126] = 13;
        pixel_data[180][127] = 13;
        pixel_data[180][128] = 13;
        pixel_data[180][129] = 13;
        pixel_data[180][130] = 13;
        pixel_data[180][131] = 13;
        pixel_data[180][132] = 13;
        pixel_data[180][133] = 13;
        pixel_data[180][134] = 13;
        pixel_data[180][135] = 13;
        pixel_data[180][136] = 10;
        pixel_data[180][137] = 5;
        pixel_data[180][138] = 1;
        pixel_data[180][139] = 1;
        pixel_data[180][140] = 1;
        pixel_data[180][141] = 1;
        pixel_data[180][142] = 1;
        pixel_data[180][143] = 1;
        pixel_data[180][144] = 1;
        pixel_data[180][145] = 1;
        pixel_data[180][146] = 1;
        pixel_data[180][147] = 1;
        pixel_data[180][148] = 1;
        pixel_data[180][149] = 1;
        pixel_data[180][150] = 1;
        pixel_data[180][151] = 1;
        pixel_data[180][152] = 1;
        pixel_data[180][153] = 1;
        pixel_data[180][154] = 1;
        pixel_data[180][155] = 1;
        pixel_data[180][156] = 1;
        pixel_data[180][157] = 1;
        pixel_data[180][158] = 1;
        pixel_data[180][159] = 1;
        pixel_data[180][160] = 1;
        pixel_data[180][161] = 1;
        pixel_data[180][162] = 1;
        pixel_data[180][163] = 1;
        pixel_data[180][164] = 1;
        pixel_data[180][165] = 1;
        pixel_data[180][166] = 1;
        pixel_data[180][167] = 1;
        pixel_data[180][168] = 1;
        pixel_data[180][169] = 1;
        pixel_data[180][170] = 1;
        pixel_data[180][171] = 1;
        pixel_data[180][172] = 1;
        pixel_data[180][173] = 1;
        pixel_data[180][174] = 1;
        pixel_data[180][175] = 1;
        pixel_data[180][176] = 1;
        pixel_data[180][177] = 1;
        pixel_data[180][178] = 1;
        pixel_data[180][179] = 1;
        pixel_data[180][180] = 1;
        pixel_data[180][181] = 1;
        pixel_data[180][182] = 1;
        pixel_data[180][183] = 1;
        pixel_data[180][184] = 1;
        pixel_data[180][185] = 1;
        pixel_data[180][186] = 1;
        pixel_data[180][187] = 6;
        pixel_data[180][188] = 9;
        pixel_data[180][189] = 11;
        pixel_data[180][190] = 11;
        pixel_data[180][191] = 0;
        pixel_data[180][192] = 0;
        pixel_data[180][193] = 0;
        pixel_data[180][194] = 0;
        pixel_data[180][195] = 0;
        pixel_data[180][196] = 0;
        pixel_data[180][197] = 0;
        pixel_data[180][198] = 0;
        pixel_data[180][199] = 0; // y=180
        pixel_data[181][0] = 0;
        pixel_data[181][1] = 0;
        pixel_data[181][2] = 0;
        pixel_data[181][3] = 0;
        pixel_data[181][4] = 11;
        pixel_data[181][5] = 11;
        pixel_data[181][6] = 9;
        pixel_data[181][7] = 6;
        pixel_data[181][8] = 1;
        pixel_data[181][9] = 1;
        pixel_data[181][10] = 1;
        pixel_data[181][11] = 1;
        pixel_data[181][12] = 2;
        pixel_data[181][13] = 4;
        pixel_data[181][14] = 4;
        pixel_data[181][15] = 1;
        pixel_data[181][16] = 1;
        pixel_data[181][17] = 1;
        pixel_data[181][18] = 1;
        pixel_data[181][19] = 1;
        pixel_data[181][20] = 1;
        pixel_data[181][21] = 1;
        pixel_data[181][22] = 1;
        pixel_data[181][23] = 1;
        pixel_data[181][24] = 1;
        pixel_data[181][25] = 1;
        pixel_data[181][26] = 1;
        pixel_data[181][27] = 1;
        pixel_data[181][28] = 1;
        pixel_data[181][29] = 1;
        pixel_data[181][30] = 1;
        pixel_data[181][31] = 1;
        pixel_data[181][32] = 1;
        pixel_data[181][33] = 1;
        pixel_data[181][34] = 1;
        pixel_data[181][35] = 1;
        pixel_data[181][36] = 1;
        pixel_data[181][37] = 1;
        pixel_data[181][38] = 1;
        pixel_data[181][39] = 1;
        pixel_data[181][40] = 1;
        pixel_data[181][41] = 1;
        pixel_data[181][42] = 1;
        pixel_data[181][43] = 1;
        pixel_data[181][44] = 1;
        pixel_data[181][45] = 1;
        pixel_data[181][46] = 1;
        pixel_data[181][47] = 1;
        pixel_data[181][48] = 1;
        pixel_data[181][49] = 1;
        pixel_data[181][50] = 1;
        pixel_data[181][51] = 1;
        pixel_data[181][52] = 1;
        pixel_data[181][53] = 1;
        pixel_data[181][54] = 1;
        pixel_data[181][55] = 1;
        pixel_data[181][56] = 1;
        pixel_data[181][57] = 1;
        pixel_data[181][58] = 1;
        pixel_data[181][59] = 1;
        pixel_data[181][60] = 1;
        pixel_data[181][61] = 1;
        pixel_data[181][62] = 1;
        pixel_data[181][63] = 1;
        pixel_data[181][64] = 1;
        pixel_data[181][65] = 1;
        pixel_data[181][66] = 1;
        pixel_data[181][67] = 1;
        pixel_data[181][68] = 1;
        pixel_data[181][69] = 1;
        pixel_data[181][70] = 1;
        pixel_data[181][71] = 1;
        pixel_data[181][72] = 1;
        pixel_data[181][73] = 1;
        pixel_data[181][74] = 1;
        pixel_data[181][75] = 1;
        pixel_data[181][76] = 1;
        pixel_data[181][77] = 1;
        pixel_data[181][78] = 1;
        pixel_data[181][79] = 1;
        pixel_data[181][80] = 1;
        pixel_data[181][81] = 1;
        pixel_data[181][82] = 1;
        pixel_data[181][83] = 1;
        pixel_data[181][84] = 1;
        pixel_data[181][85] = 1;
        pixel_data[181][86] = 1;
        pixel_data[181][87] = 1;
        pixel_data[181][88] = 1;
        pixel_data[181][89] = 1;
        pixel_data[181][90] = 1;
        pixel_data[181][91] = 1;
        pixel_data[181][92] = 1;
        pixel_data[181][93] = 1;
        pixel_data[181][94] = 1;
        pixel_data[181][95] = 1;
        pixel_data[181][96] = 1;
        pixel_data[181][97] = 1;
        pixel_data[181][98] = 1;
        pixel_data[181][99] = 1;
        pixel_data[181][100] = 1;
        pixel_data[181][101] = 1;
        pixel_data[181][102] = 1;
        pixel_data[181][103] = 1;
        pixel_data[181][104] = 1;
        pixel_data[181][105] = 1;
        pixel_data[181][106] = 1;
        pixel_data[181][107] = 1;
        pixel_data[181][108] = 1;
        pixel_data[181][109] = 1;
        pixel_data[181][110] = 1;
        pixel_data[181][111] = 1;
        pixel_data[181][112] = 1;
        pixel_data[181][113] = 7;
        pixel_data[181][114] = 10;
        pixel_data[181][115] = 13;
        pixel_data[181][116] = 13;
        pixel_data[181][117] = 13;
        pixel_data[181][118] = 13;
        pixel_data[181][119] = 13;
        pixel_data[181][120] = 13;
        pixel_data[181][121] = 13;
        pixel_data[181][122] = 13;
        pixel_data[181][123] = 13;
        pixel_data[181][124] = 13;
        pixel_data[181][125] = 13;
        pixel_data[181][126] = 13;
        pixel_data[181][127] = 13;
        pixel_data[181][128] = 13;
        pixel_data[181][129] = 13;
        pixel_data[181][130] = 13;
        pixel_data[181][131] = 13;
        pixel_data[181][132] = 13;
        pixel_data[181][133] = 13;
        pixel_data[181][134] = 13;
        pixel_data[181][135] = 10;
        pixel_data[181][136] = 7;
        pixel_data[181][137] = 1;
        pixel_data[181][138] = 1;
        pixel_data[181][139] = 1;
        pixel_data[181][140] = 1;
        pixel_data[181][141] = 1;
        pixel_data[181][142] = 1;
        pixel_data[181][143] = 1;
        pixel_data[181][144] = 1;
        pixel_data[181][145] = 1;
        pixel_data[181][146] = 1;
        pixel_data[181][147] = 1;
        pixel_data[181][148] = 1;
        pixel_data[181][149] = 1;
        pixel_data[181][150] = 1;
        pixel_data[181][151] = 1;
        pixel_data[181][152] = 1;
        pixel_data[181][153] = 1;
        pixel_data[181][154] = 1;
        pixel_data[181][155] = 1;
        pixel_data[181][156] = 1;
        pixel_data[181][157] = 1;
        pixel_data[181][158] = 1;
        pixel_data[181][159] = 1;
        pixel_data[181][160] = 1;
        pixel_data[181][161] = 1;
        pixel_data[181][162] = 1;
        pixel_data[181][163] = 1;
        pixel_data[181][164] = 1;
        pixel_data[181][165] = 1;
        pixel_data[181][166] = 1;
        pixel_data[181][167] = 1;
        pixel_data[181][168] = 1;
        pixel_data[181][169] = 1;
        pixel_data[181][170] = 1;
        pixel_data[181][171] = 1;
        pixel_data[181][172] = 1;
        pixel_data[181][173] = 1;
        pixel_data[181][174] = 1;
        pixel_data[181][175] = 1;
        pixel_data[181][176] = 1;
        pixel_data[181][177] = 1;
        pixel_data[181][178] = 1;
        pixel_data[181][179] = 1;
        pixel_data[181][180] = 1;
        pixel_data[181][181] = 1;
        pixel_data[181][182] = 1;
        pixel_data[181][183] = 1;
        pixel_data[181][184] = 1;
        pixel_data[181][185] = 1;
        pixel_data[181][186] = 1;
        pixel_data[181][187] = 5;
        pixel_data[181][188] = 8;
        pixel_data[181][189] = 11;
        pixel_data[181][190] = 11;
        pixel_data[181][191] = 0;
        pixel_data[181][192] = 0;
        pixel_data[181][193] = 0;
        pixel_data[181][194] = 0;
        pixel_data[181][195] = 0;
        pixel_data[181][196] = 0;
        pixel_data[181][197] = 0;
        pixel_data[181][198] = 0;
        pixel_data[181][199] = 0; // y=181
        pixel_data[182][0] = 0;
        pixel_data[182][1] = 0;
        pixel_data[182][2] = 0;
        pixel_data[182][3] = 0;
        pixel_data[182][4] = 11;
        pixel_data[182][5] = 11;
        pixel_data[182][6] = 9;
        pixel_data[182][7] = 6;
        pixel_data[182][8] = 1;
        pixel_data[182][9] = 1;
        pixel_data[182][10] = 1;
        pixel_data[182][11] = 1;
        pixel_data[182][12] = 2;
        pixel_data[182][13] = 4;
        pixel_data[182][14] = 4;
        pixel_data[182][15] = 1;
        pixel_data[182][16] = 1;
        pixel_data[182][17] = 1;
        pixel_data[182][18] = 1;
        pixel_data[182][19] = 1;
        pixel_data[182][20] = 1;
        pixel_data[182][21] = 1;
        pixel_data[182][22] = 1;
        pixel_data[182][23] = 1;
        pixel_data[182][24] = 1;
        pixel_data[182][25] = 1;
        pixel_data[182][26] = 1;
        pixel_data[182][27] = 1;
        pixel_data[182][28] = 1;
        pixel_data[182][29] = 1;
        pixel_data[182][30] = 1;
        pixel_data[182][31] = 1;
        pixel_data[182][32] = 1;
        pixel_data[182][33] = 1;
        pixel_data[182][34] = 1;
        pixel_data[182][35] = 1;
        pixel_data[182][36] = 1;
        pixel_data[182][37] = 1;
        pixel_data[182][38] = 1;
        pixel_data[182][39] = 1;
        pixel_data[182][40] = 1;
        pixel_data[182][41] = 1;
        pixel_data[182][42] = 1;
        pixel_data[182][43] = 1;
        pixel_data[182][44] = 1;
        pixel_data[182][45] = 1;
        pixel_data[182][46] = 1;
        pixel_data[182][47] = 1;
        pixel_data[182][48] = 1;
        pixel_data[182][49] = 1;
        pixel_data[182][50] = 1;
        pixel_data[182][51] = 1;
        pixel_data[182][52] = 1;
        pixel_data[182][53] = 1;
        pixel_data[182][54] = 1;
        pixel_data[182][55] = 1;
        pixel_data[182][56] = 1;
        pixel_data[182][57] = 1;
        pixel_data[182][58] = 1;
        pixel_data[182][59] = 1;
        pixel_data[182][60] = 1;
        pixel_data[182][61] = 1;
        pixel_data[182][62] = 1;
        pixel_data[182][63] = 1;
        pixel_data[182][64] = 1;
        pixel_data[182][65] = 1;
        pixel_data[182][66] = 1;
        pixel_data[182][67] = 1;
        pixel_data[182][68] = 1;
        pixel_data[182][69] = 1;
        pixel_data[182][70] = 1;
        pixel_data[182][71] = 1;
        pixel_data[182][72] = 1;
        pixel_data[182][73] = 1;
        pixel_data[182][74] = 1;
        pixel_data[182][75] = 1;
        pixel_data[182][76] = 1;
        pixel_data[182][77] = 1;
        pixel_data[182][78] = 1;
        pixel_data[182][79] = 1;
        pixel_data[182][80] = 1;
        pixel_data[182][81] = 1;
        pixel_data[182][82] = 1;
        pixel_data[182][83] = 1;
        pixel_data[182][84] = 1;
        pixel_data[182][85] = 1;
        pixel_data[182][86] = 1;
        pixel_data[182][87] = 1;
        pixel_data[182][88] = 1;
        pixel_data[182][89] = 1;
        pixel_data[182][90] = 1;
        pixel_data[182][91] = 1;
        pixel_data[182][92] = 1;
        pixel_data[182][93] = 1;
        pixel_data[182][94] = 1;
        pixel_data[182][95] = 1;
        pixel_data[182][96] = 1;
        pixel_data[182][97] = 1;
        pixel_data[182][98] = 1;
        pixel_data[182][99] = 1;
        pixel_data[182][100] = 1;
        pixel_data[182][101] = 1;
        pixel_data[182][102] = 1;
        pixel_data[182][103] = 1;
        pixel_data[182][104] = 1;
        pixel_data[182][105] = 1;
        pixel_data[182][106] = 1;
        pixel_data[182][107] = 1;
        pixel_data[182][108] = 1;
        pixel_data[182][109] = 1;
        pixel_data[182][110] = 1;
        pixel_data[182][111] = 1;
        pixel_data[182][112] = 1;
        pixel_data[182][113] = 1;
        pixel_data[182][114] = 5;
        pixel_data[182][115] = 8;
        pixel_data[182][116] = 12;
        pixel_data[182][117] = 13;
        pixel_data[182][118] = 13;
        pixel_data[182][119] = 13;
        pixel_data[182][120] = 13;
        pixel_data[182][121] = 13;
        pixel_data[182][122] = 13;
        pixel_data[182][123] = 13;
        pixel_data[182][124] = 13;
        pixel_data[182][125] = 13;
        pixel_data[182][126] = 13;
        pixel_data[182][127] = 13;
        pixel_data[182][128] = 13;
        pixel_data[182][129] = 13;
        pixel_data[182][130] = 13;
        pixel_data[182][131] = 13;
        pixel_data[182][132] = 13;
        pixel_data[182][133] = 13;
        pixel_data[182][134] = 10;
        pixel_data[182][135] = 5;
        pixel_data[182][136] = 1;
        pixel_data[182][137] = 1;
        pixel_data[182][138] = 1;
        pixel_data[182][139] = 1;
        pixel_data[182][140] = 1;
        pixel_data[182][141] = 1;
        pixel_data[182][142] = 1;
        pixel_data[182][143] = 1;
        pixel_data[182][144] = 1;
        pixel_data[182][145] = 1;
        pixel_data[182][146] = 1;
        pixel_data[182][147] = 1;
        pixel_data[182][148] = 1;
        pixel_data[182][149] = 1;
        pixel_data[182][150] = 1;
        pixel_data[182][151] = 1;
        pixel_data[182][152] = 1;
        pixel_data[182][153] = 1;
        pixel_data[182][154] = 1;
        pixel_data[182][155] = 1;
        pixel_data[182][156] = 1;
        pixel_data[182][157] = 1;
        pixel_data[182][158] = 1;
        pixel_data[182][159] = 1;
        pixel_data[182][160] = 1;
        pixel_data[182][161] = 1;
        pixel_data[182][162] = 1;
        pixel_data[182][163] = 1;
        pixel_data[182][164] = 1;
        pixel_data[182][165] = 1;
        pixel_data[182][166] = 1;
        pixel_data[182][167] = 1;
        pixel_data[182][168] = 1;
        pixel_data[182][169] = 1;
        pixel_data[182][170] = 1;
        pixel_data[182][171] = 1;
        pixel_data[182][172] = 1;
        pixel_data[182][173] = 1;
        pixel_data[182][174] = 1;
        pixel_data[182][175] = 1;
        pixel_data[182][176] = 1;
        pixel_data[182][177] = 1;
        pixel_data[182][178] = 1;
        pixel_data[182][179] = 1;
        pixel_data[182][180] = 1;
        pixel_data[182][181] = 1;
        pixel_data[182][182] = 1;
        pixel_data[182][183] = 1;
        pixel_data[182][184] = 1;
        pixel_data[182][185] = 1;
        pixel_data[182][186] = 1;
        pixel_data[182][187] = 1;
        pixel_data[182][188] = 6;
        pixel_data[182][189] = 8;
        pixel_data[182][190] = 11;
        pixel_data[182][191] = 11;
        pixel_data[182][192] = 0;
        pixel_data[182][193] = 0;
        pixel_data[182][194] = 0;
        pixel_data[182][195] = 0;
        pixel_data[182][196] = 0;
        pixel_data[182][197] = 0;
        pixel_data[182][198] = 0;
        pixel_data[182][199] = 0; // y=182
        pixel_data[183][0] = 0;
        pixel_data[183][1] = 0;
        pixel_data[183][2] = 0;
        pixel_data[183][3] = 0;
        pixel_data[183][4] = 11;
        pixel_data[183][5] = 11;
        pixel_data[183][6] = 8;
        pixel_data[183][7] = 4;
        pixel_data[183][8] = 1;
        pixel_data[183][9] = 1;
        pixel_data[183][10] = 1;
        pixel_data[183][11] = 1;
        pixel_data[183][12] = 2;
        pixel_data[183][13] = 4;
        pixel_data[183][14] = 4;
        pixel_data[183][15] = 1;
        pixel_data[183][16] = 1;
        pixel_data[183][17] = 1;
        pixel_data[183][18] = 1;
        pixel_data[183][19] = 1;
        pixel_data[183][20] = 1;
        pixel_data[183][21] = 1;
        pixel_data[183][22] = 1;
        pixel_data[183][23] = 1;
        pixel_data[183][24] = 1;
        pixel_data[183][25] = 1;
        pixel_data[183][26] = 1;
        pixel_data[183][27] = 1;
        pixel_data[183][28] = 1;
        pixel_data[183][29] = 1;
        pixel_data[183][30] = 1;
        pixel_data[183][31] = 1;
        pixel_data[183][32] = 1;
        pixel_data[183][33] = 1;
        pixel_data[183][34] = 1;
        pixel_data[183][35] = 1;
        pixel_data[183][36] = 1;
        pixel_data[183][37] = 1;
        pixel_data[183][38] = 1;
        pixel_data[183][39] = 1;
        pixel_data[183][40] = 1;
        pixel_data[183][41] = 1;
        pixel_data[183][42] = 1;
        pixel_data[183][43] = 1;
        pixel_data[183][44] = 1;
        pixel_data[183][45] = 1;
        pixel_data[183][46] = 1;
        pixel_data[183][47] = 1;
        pixel_data[183][48] = 1;
        pixel_data[183][49] = 1;
        pixel_data[183][50] = 1;
        pixel_data[183][51] = 1;
        pixel_data[183][52] = 1;
        pixel_data[183][53] = 1;
        pixel_data[183][54] = 1;
        pixel_data[183][55] = 1;
        pixel_data[183][56] = 1;
        pixel_data[183][57] = 1;
        pixel_data[183][58] = 1;
        pixel_data[183][59] = 1;
        pixel_data[183][60] = 1;
        pixel_data[183][61] = 1;
        pixel_data[183][62] = 1;
        pixel_data[183][63] = 1;
        pixel_data[183][64] = 1;
        pixel_data[183][65] = 1;
        pixel_data[183][66] = 1;
        pixel_data[183][67] = 1;
        pixel_data[183][68] = 1;
        pixel_data[183][69] = 1;
        pixel_data[183][70] = 1;
        pixel_data[183][71] = 1;
        pixel_data[183][72] = 1;
        pixel_data[183][73] = 1;
        pixel_data[183][74] = 1;
        pixel_data[183][75] = 1;
        pixel_data[183][76] = 1;
        pixel_data[183][77] = 1;
        pixel_data[183][78] = 1;
        pixel_data[183][79] = 1;
        pixel_data[183][80] = 1;
        pixel_data[183][81] = 1;
        pixel_data[183][82] = 1;
        pixel_data[183][83] = 1;
        pixel_data[183][84] = 1;
        pixel_data[183][85] = 1;
        pixel_data[183][86] = 1;
        pixel_data[183][87] = 1;
        pixel_data[183][88] = 1;
        pixel_data[183][89] = 1;
        pixel_data[183][90] = 1;
        pixel_data[183][91] = 1;
        pixel_data[183][92] = 1;
        pixel_data[183][93] = 1;
        pixel_data[183][94] = 1;
        pixel_data[183][95] = 1;
        pixel_data[183][96] = 1;
        pixel_data[183][97] = 1;
        pixel_data[183][98] = 1;
        pixel_data[183][99] = 1;
        pixel_data[183][100] = 1;
        pixel_data[183][101] = 1;
        pixel_data[183][102] = 1;
        pixel_data[183][103] = 1;
        pixel_data[183][104] = 1;
        pixel_data[183][105] = 1;
        pixel_data[183][106] = 1;
        pixel_data[183][107] = 1;
        pixel_data[183][108] = 1;
        pixel_data[183][109] = 1;
        pixel_data[183][110] = 1;
        pixel_data[183][111] = 1;
        pixel_data[183][112] = 1;
        pixel_data[183][113] = 1;
        pixel_data[183][114] = 1;
        pixel_data[183][115] = 1;
        pixel_data[183][116] = 5;
        pixel_data[183][117] = 9;
        pixel_data[183][118] = 12;
        pixel_data[183][119] = 13;
        pixel_data[183][120] = 13;
        pixel_data[183][121] = 13;
        pixel_data[183][122] = 13;
        pixel_data[183][123] = 13;
        pixel_data[183][124] = 13;
        pixel_data[183][125] = 13;
        pixel_data[183][126] = 13;
        pixel_data[183][127] = 13;
        pixel_data[183][128] = 13;
        pixel_data[183][129] = 13;
        pixel_data[183][130] = 13;
        pixel_data[183][131] = 13;
        pixel_data[183][132] = 12;
        pixel_data[183][133] = 7;
        pixel_data[183][134] = 1;
        pixel_data[183][135] = 1;
        pixel_data[183][136] = 1;
        pixel_data[183][137] = 1;
        pixel_data[183][138] = 1;
        pixel_data[183][139] = 1;
        pixel_data[183][140] = 1;
        pixel_data[183][141] = 1;
        pixel_data[183][142] = 1;
        pixel_data[183][143] = 1;
        pixel_data[183][144] = 1;
        pixel_data[183][145] = 1;
        pixel_data[183][146] = 1;
        pixel_data[183][147] = 1;
        pixel_data[183][148] = 1;
        pixel_data[183][149] = 1;
        pixel_data[183][150] = 1;
        pixel_data[183][151] = 1;
        pixel_data[183][152] = 1;
        pixel_data[183][153] = 1;
        pixel_data[183][154] = 1;
        pixel_data[183][155] = 1;
        pixel_data[183][156] = 1;
        pixel_data[183][157] = 1;
        pixel_data[183][158] = 1;
        pixel_data[183][159] = 1;
        pixel_data[183][160] = 1;
        pixel_data[183][161] = 1;
        pixel_data[183][162] = 1;
        pixel_data[183][163] = 1;
        pixel_data[183][164] = 1;
        pixel_data[183][165] = 1;
        pixel_data[183][166] = 1;
        pixel_data[183][167] = 1;
        pixel_data[183][168] = 1;
        pixel_data[183][169] = 1;
        pixel_data[183][170] = 1;
        pixel_data[183][171] = 1;
        pixel_data[183][172] = 1;
        pixel_data[183][173] = 1;
        pixel_data[183][174] = 1;
        pixel_data[183][175] = 1;
        pixel_data[183][176] = 1;
        pixel_data[183][177] = 1;
        pixel_data[183][178] = 1;
        pixel_data[183][179] = 1;
        pixel_data[183][180] = 1;
        pixel_data[183][181] = 1;
        pixel_data[183][182] = 1;
        pixel_data[183][183] = 1;
        pixel_data[183][184] = 1;
        pixel_data[183][185] = 1;
        pixel_data[183][186] = 1;
        pixel_data[183][187] = 1;
        pixel_data[183][188] = 4;
        pixel_data[183][189] = 7;
        pixel_data[183][190] = 11;
        pixel_data[183][191] = 11;
        pixel_data[183][192] = 0;
        pixel_data[183][193] = 0;
        pixel_data[183][194] = 0;
        pixel_data[183][195] = 0;
        pixel_data[183][196] = 0;
        pixel_data[183][197] = 0;
        pixel_data[183][198] = 0;
        pixel_data[183][199] = 0; // y=183
        pixel_data[184][0] = 0;
        pixel_data[184][1] = 0;
        pixel_data[184][2] = 0;
        pixel_data[184][3] = 0;
        pixel_data[184][4] = 11;
        pixel_data[184][5] = 11;
        pixel_data[184][6] = 8;
        pixel_data[184][7] = 4;
        pixel_data[184][8] = 1;
        pixel_data[184][9] = 1;
        pixel_data[184][10] = 1;
        pixel_data[184][11] = 1;
        pixel_data[184][12] = 2;
        pixel_data[184][13] = 4;
        pixel_data[184][14] = 4;
        pixel_data[184][15] = 1;
        pixel_data[184][16] = 1;
        pixel_data[184][17] = 1;
        pixel_data[184][18] = 1;
        pixel_data[184][19] = 1;
        pixel_data[184][20] = 1;
        pixel_data[184][21] = 1;
        pixel_data[184][22] = 1;
        pixel_data[184][23] = 1;
        pixel_data[184][24] = 1;
        pixel_data[184][25] = 1;
        pixel_data[184][26] = 1;
        pixel_data[184][27] = 1;
        pixel_data[184][28] = 1;
        pixel_data[184][29] = 1;
        pixel_data[184][30] = 1;
        pixel_data[184][31] = 1;
        pixel_data[184][32] = 1;
        pixel_data[184][33] = 1;
        pixel_data[184][34] = 1;
        pixel_data[184][35] = 1;
        pixel_data[184][36] = 1;
        pixel_data[184][37] = 1;
        pixel_data[184][38] = 1;
        pixel_data[184][39] = 1;
        pixel_data[184][40] = 1;
        pixel_data[184][41] = 1;
        pixel_data[184][42] = 1;
        pixel_data[184][43] = 1;
        pixel_data[184][44] = 1;
        pixel_data[184][45] = 1;
        pixel_data[184][46] = 1;
        pixel_data[184][47] = 1;
        pixel_data[184][48] = 1;
        pixel_data[184][49] = 1;
        pixel_data[184][50] = 1;
        pixel_data[184][51] = 1;
        pixel_data[184][52] = 1;
        pixel_data[184][53] = 1;
        pixel_data[184][54] = 1;
        pixel_data[184][55] = 1;
        pixel_data[184][56] = 1;
        pixel_data[184][57] = 1;
        pixel_data[184][58] = 1;
        pixel_data[184][59] = 1;
        pixel_data[184][60] = 1;
        pixel_data[184][61] = 1;
        pixel_data[184][62] = 1;
        pixel_data[184][63] = 1;
        pixel_data[184][64] = 1;
        pixel_data[184][65] = 1;
        pixel_data[184][66] = 1;
        pixel_data[184][67] = 1;
        pixel_data[184][68] = 1;
        pixel_data[184][69] = 1;
        pixel_data[184][70] = 1;
        pixel_data[184][71] = 1;
        pixel_data[184][72] = 1;
        pixel_data[184][73] = 1;
        pixel_data[184][74] = 1;
        pixel_data[184][75] = 1;
        pixel_data[184][76] = 1;
        pixel_data[184][77] = 1;
        pixel_data[184][78] = 1;
        pixel_data[184][79] = 1;
        pixel_data[184][80] = 1;
        pixel_data[184][81] = 1;
        pixel_data[184][82] = 1;
        pixel_data[184][83] = 1;
        pixel_data[184][84] = 1;
        pixel_data[184][85] = 1;
        pixel_data[184][86] = 1;
        pixel_data[184][87] = 1;
        pixel_data[184][88] = 1;
        pixel_data[184][89] = 1;
        pixel_data[184][90] = 1;
        pixel_data[184][91] = 1;
        pixel_data[184][92] = 1;
        pixel_data[184][93] = 1;
        pixel_data[184][94] = 1;
        pixel_data[184][95] = 1;
        pixel_data[184][96] = 1;
        pixel_data[184][97] = 1;
        pixel_data[184][98] = 1;
        pixel_data[184][99] = 1;
        pixel_data[184][100] = 1;
        pixel_data[184][101] = 1;
        pixel_data[184][102] = 1;
        pixel_data[184][103] = 1;
        pixel_data[184][104] = 1;
        pixel_data[184][105] = 1;
        pixel_data[184][106] = 1;
        pixel_data[184][107] = 1;
        pixel_data[184][108] = 1;
        pixel_data[184][109] = 1;
        pixel_data[184][110] = 1;
        pixel_data[184][111] = 1;
        pixel_data[184][112] = 1;
        pixel_data[184][113] = 1;
        pixel_data[184][114] = 1;
        pixel_data[184][115] = 1;
        pixel_data[184][116] = 1;
        pixel_data[184][117] = 1;
        pixel_data[184][118] = 1;
        pixel_data[184][119] = 6;
        pixel_data[184][120] = 9;
        pixel_data[184][121] = 12;
        pixel_data[184][122] = 13;
        pixel_data[184][123] = 13;
        pixel_data[184][124] = 13;
        pixel_data[184][125] = 13;
        pixel_data[184][126] = 13;
        pixel_data[184][127] = 13;
        pixel_data[184][128] = 13;
        pixel_data[184][129] = 13;
        pixel_data[184][130] = 12;
        pixel_data[184][131] = 9;
        pixel_data[184][132] = 4;
        pixel_data[184][133] = 1;
        pixel_data[184][134] = 1;
        pixel_data[184][135] = 1;
        pixel_data[184][136] = 1;
        pixel_data[184][137] = 1;
        pixel_data[184][138] = 1;
        pixel_data[184][139] = 1;
        pixel_data[184][140] = 1;
        pixel_data[184][141] = 1;
        pixel_data[184][142] = 1;
        pixel_data[184][143] = 1;
        pixel_data[184][144] = 1;
        pixel_data[184][145] = 1;
        pixel_data[184][146] = 1;
        pixel_data[184][147] = 1;
        pixel_data[184][148] = 1;
        pixel_data[184][149] = 1;
        pixel_data[184][150] = 1;
        pixel_data[184][151] = 1;
        pixel_data[184][152] = 1;
        pixel_data[184][153] = 1;
        pixel_data[184][154] = 1;
        pixel_data[184][155] = 1;
        pixel_data[184][156] = 1;
        pixel_data[184][157] = 1;
        pixel_data[184][158] = 1;
        pixel_data[184][159] = 1;
        pixel_data[184][160] = 1;
        pixel_data[184][161] = 1;
        pixel_data[184][162] = 1;
        pixel_data[184][163] = 1;
        pixel_data[184][164] = 1;
        pixel_data[184][165] = 1;
        pixel_data[184][166] = 1;
        pixel_data[184][167] = 1;
        pixel_data[184][168] = 1;
        pixel_data[184][169] = 1;
        pixel_data[184][170] = 1;
        pixel_data[184][171] = 1;
        pixel_data[184][172] = 1;
        pixel_data[184][173] = 1;
        pixel_data[184][174] = 1;
        pixel_data[184][175] = 1;
        pixel_data[184][176] = 1;
        pixel_data[184][177] = 1;
        pixel_data[184][178] = 1;
        pixel_data[184][179] = 1;
        pixel_data[184][180] = 1;
        pixel_data[184][181] = 1;
        pixel_data[184][182] = 1;
        pixel_data[184][183] = 1;
        pixel_data[184][184] = 1;
        pixel_data[184][185] = 1;
        pixel_data[184][186] = 1;
        pixel_data[184][187] = 1;
        pixel_data[184][188] = 1;
        pixel_data[184][189] = 6;
        pixel_data[184][190] = 9;
        pixel_data[184][191] = 11;
        pixel_data[184][192] = 11;
        pixel_data[184][193] = 0;
        pixel_data[184][194] = 0;
        pixel_data[184][195] = 0;
        pixel_data[184][196] = 0;
        pixel_data[184][197] = 0;
        pixel_data[184][198] = 0;
        pixel_data[184][199] = 0; // y=184
        pixel_data[185][0] = 0;
        pixel_data[185][1] = 0;
        pixel_data[185][2] = 0;
        pixel_data[185][3] = 10;
        pixel_data[185][4] = 11;
        pixel_data[185][5] = 11;
        pixel_data[185][6] = 7;
        pixel_data[185][7] = 1;
        pixel_data[185][8] = 1;
        pixel_data[185][9] = 1;
        pixel_data[185][10] = 1;
        pixel_data[185][11] = 1;
        pixel_data[185][12] = 1;
        pixel_data[185][13] = 4;
        pixel_data[185][14] = 4;
        pixel_data[185][15] = 2;
        pixel_data[185][16] = 1;
        pixel_data[185][17] = 1;
        pixel_data[185][18] = 1;
        pixel_data[185][19] = 1;
        pixel_data[185][20] = 1;
        pixel_data[185][21] = 1;
        pixel_data[185][22] = 1;
        pixel_data[185][23] = 1;
        pixel_data[185][24] = 1;
        pixel_data[185][25] = 1;
        pixel_data[185][26] = 1;
        pixel_data[185][27] = 1;
        pixel_data[185][28] = 1;
        pixel_data[185][29] = 1;
        pixel_data[185][30] = 1;
        pixel_data[185][31] = 1;
        pixel_data[185][32] = 1;
        pixel_data[185][33] = 1;
        pixel_data[185][34] = 1;
        pixel_data[185][35] = 1;
        pixel_data[185][36] = 1;
        pixel_data[185][37] = 1;
        pixel_data[185][38] = 1;
        pixel_data[185][39] = 1;
        pixel_data[185][40] = 1;
        pixel_data[185][41] = 1;
        pixel_data[185][42] = 1;
        pixel_data[185][43] = 1;
        pixel_data[185][44] = 1;
        pixel_data[185][45] = 1;
        pixel_data[185][46] = 1;
        pixel_data[185][47] = 1;
        pixel_data[185][48] = 1;
        pixel_data[185][49] = 1;
        pixel_data[185][50] = 1;
        pixel_data[185][51] = 1;
        pixel_data[185][52] = 1;
        pixel_data[185][53] = 1;
        pixel_data[185][54] = 1;
        pixel_data[185][55] = 1;
        pixel_data[185][56] = 1;
        pixel_data[185][57] = 1;
        pixel_data[185][58] = 1;
        pixel_data[185][59] = 1;
        pixel_data[185][60] = 1;
        pixel_data[185][61] = 1;
        pixel_data[185][62] = 1;
        pixel_data[185][63] = 1;
        pixel_data[185][64] = 1;
        pixel_data[185][65] = 1;
        pixel_data[185][66] = 1;
        pixel_data[185][67] = 1;
        pixel_data[185][68] = 1;
        pixel_data[185][69] = 1;
        pixel_data[185][70] = 1;
        pixel_data[185][71] = 1;
        pixel_data[185][72] = 1;
        pixel_data[185][73] = 1;
        pixel_data[185][74] = 1;
        pixel_data[185][75] = 1;
        pixel_data[185][76] = 1;
        pixel_data[185][77] = 1;
        pixel_data[185][78] = 1;
        pixel_data[185][79] = 1;
        pixel_data[185][80] = 1;
        pixel_data[185][81] = 1;
        pixel_data[185][82] = 1;
        pixel_data[185][83] = 1;
        pixel_data[185][84] = 1;
        pixel_data[185][85] = 1;
        pixel_data[185][86] = 1;
        pixel_data[185][87] = 1;
        pixel_data[185][88] = 1;
        pixel_data[185][89] = 1;
        pixel_data[185][90] = 1;
        pixel_data[185][91] = 1;
        pixel_data[185][92] = 1;
        pixel_data[185][93] = 1;
        pixel_data[185][94] = 1;
        pixel_data[185][95] = 1;
        pixel_data[185][96] = 1;
        pixel_data[185][97] = 1;
        pixel_data[185][98] = 1;
        pixel_data[185][99] = 1;
        pixel_data[185][100] = 1;
        pixel_data[185][101] = 1;
        pixel_data[185][102] = 1;
        pixel_data[185][103] = 1;
        pixel_data[185][104] = 1;
        pixel_data[185][105] = 1;
        pixel_data[185][106] = 1;
        pixel_data[185][107] = 1;
        pixel_data[185][108] = 1;
        pixel_data[185][109] = 1;
        pixel_data[185][110] = 1;
        pixel_data[185][111] = 1;
        pixel_data[185][112] = 1;
        pixel_data[185][113] = 1;
        pixel_data[185][114] = 1;
        pixel_data[185][115] = 1;
        pixel_data[185][116] = 1;
        pixel_data[185][117] = 1;
        pixel_data[185][118] = 1;
        pixel_data[185][119] = 1;
        pixel_data[185][120] = 1;
        pixel_data[185][121] = 1;
        pixel_data[185][122] = 1;
        pixel_data[185][123] = 1;
        pixel_data[185][124] = 1;
        pixel_data[185][125] = 1;
        pixel_data[185][126] = 4;
        pixel_data[185][127] = 4;
        pixel_data[185][128] = 1;
        pixel_data[185][129] = 1;
        pixel_data[185][130] = 1;
        pixel_data[185][131] = 1;
        pixel_data[185][132] = 1;
        pixel_data[185][133] = 1;
        pixel_data[185][134] = 1;
        pixel_data[185][135] = 1;
        pixel_data[185][136] = 1;
        pixel_data[185][137] = 1;
        pixel_data[185][138] = 1;
        pixel_data[185][139] = 1;
        pixel_data[185][140] = 1;
        pixel_data[185][141] = 1;
        pixel_data[185][142] = 1;
        pixel_data[185][143] = 1;
        pixel_data[185][144] = 1;
        pixel_data[185][145] = 1;
        pixel_data[185][146] = 1;
        pixel_data[185][147] = 1;
        pixel_data[185][148] = 1;
        pixel_data[185][149] = 1;
        pixel_data[185][150] = 1;
        pixel_data[185][151] = 1;
        pixel_data[185][152] = 1;
        pixel_data[185][153] = 1;
        pixel_data[185][154] = 1;
        pixel_data[185][155] = 1;
        pixel_data[185][156] = 1;
        pixel_data[185][157] = 1;
        pixel_data[185][158] = 1;
        pixel_data[185][159] = 1;
        pixel_data[185][160] = 1;
        pixel_data[185][161] = 1;
        pixel_data[185][162] = 1;
        pixel_data[185][163] = 1;
        pixel_data[185][164] = 1;
        pixel_data[185][165] = 1;
        pixel_data[185][166] = 1;
        pixel_data[185][167] = 1;
        pixel_data[185][168] = 1;
        pixel_data[185][169] = 1;
        pixel_data[185][170] = 1;
        pixel_data[185][171] = 1;
        pixel_data[185][172] = 1;
        pixel_data[185][173] = 1;
        pixel_data[185][174] = 1;
        pixel_data[185][175] = 1;
        pixel_data[185][176] = 1;
        pixel_data[185][177] = 1;
        pixel_data[185][178] = 1;
        pixel_data[185][179] = 1;
        pixel_data[185][180] = 1;
        pixel_data[185][181] = 1;
        pixel_data[185][182] = 1;
        pixel_data[185][183] = 1;
        pixel_data[185][184] = 1;
        pixel_data[185][185] = 1;
        pixel_data[185][186] = 1;
        pixel_data[185][187] = 1;
        pixel_data[185][188] = 1;
        pixel_data[185][189] = 5;
        pixel_data[185][190] = 8;
        pixel_data[185][191] = 11;
        pixel_data[185][192] = 11;
        pixel_data[185][193] = 0;
        pixel_data[185][194] = 0;
        pixel_data[185][195] = 0;
        pixel_data[185][196] = 0;
        pixel_data[185][197] = 0;
        pixel_data[185][198] = 0;
        pixel_data[185][199] = 0; // y=185
        pixel_data[186][0] = 0;
        pixel_data[186][1] = 0;
        pixel_data[186][2] = 0;
        pixel_data[186][3] = 10;
        pixel_data[186][4] = 11;
        pixel_data[186][5] = 11;
        pixel_data[186][6] = 7;
        pixel_data[186][7] = 1;
        pixel_data[186][8] = 1;
        pixel_data[186][9] = 1;
        pixel_data[186][10] = 1;
        pixel_data[186][11] = 1;
        pixel_data[186][12] = 1;
        pixel_data[186][13] = 4;
        pixel_data[186][14] = 4;
        pixel_data[186][15] = 4;
        pixel_data[186][16] = 1;
        pixel_data[186][17] = 1;
        pixel_data[186][18] = 1;
        pixel_data[186][19] = 1;
        pixel_data[186][20] = 1;
        pixel_data[186][21] = 1;
        pixel_data[186][22] = 1;
        pixel_data[186][23] = 1;
        pixel_data[186][24] = 1;
        pixel_data[186][25] = 1;
        pixel_data[186][26] = 1;
        pixel_data[186][27] = 1;
        pixel_data[186][28] = 1;
        pixel_data[186][29] = 1;
        pixel_data[186][30] = 1;
        pixel_data[186][31] = 1;
        pixel_data[186][32] = 1;
        pixel_data[186][33] = 1;
        pixel_data[186][34] = 1;
        pixel_data[186][35] = 1;
        pixel_data[186][36] = 1;
        pixel_data[186][37] = 1;
        pixel_data[186][38] = 1;
        pixel_data[186][39] = 1;
        pixel_data[186][40] = 1;
        pixel_data[186][41] = 1;
        pixel_data[186][42] = 1;
        pixel_data[186][43] = 1;
        pixel_data[186][44] = 1;
        pixel_data[186][45] = 1;
        pixel_data[186][46] = 1;
        pixel_data[186][47] = 1;
        pixel_data[186][48] = 1;
        pixel_data[186][49] = 1;
        pixel_data[186][50] = 1;
        pixel_data[186][51] = 1;
        pixel_data[186][52] = 1;
        pixel_data[186][53] = 1;
        pixel_data[186][54] = 1;
        pixel_data[186][55] = 1;
        pixel_data[186][56] = 1;
        pixel_data[186][57] = 1;
        pixel_data[186][58] = 1;
        pixel_data[186][59] = 1;
        pixel_data[186][60] = 1;
        pixel_data[186][61] = 1;
        pixel_data[186][62] = 1;
        pixel_data[186][63] = 1;
        pixel_data[186][64] = 1;
        pixel_data[186][65] = 1;
        pixel_data[186][66] = 1;
        pixel_data[186][67] = 1;
        pixel_data[186][68] = 1;
        pixel_data[186][69] = 1;
        pixel_data[186][70] = 1;
        pixel_data[186][71] = 1;
        pixel_data[186][72] = 1;
        pixel_data[186][73] = 1;
        pixel_data[186][74] = 1;
        pixel_data[186][75] = 1;
        pixel_data[186][76] = 1;
        pixel_data[186][77] = 1;
        pixel_data[186][78] = 1;
        pixel_data[186][79] = 1;
        pixel_data[186][80] = 1;
        pixel_data[186][81] = 1;
        pixel_data[186][82] = 1;
        pixel_data[186][83] = 1;
        pixel_data[186][84] = 1;
        pixel_data[186][85] = 1;
        pixel_data[186][86] = 1;
        pixel_data[186][87] = 1;
        pixel_data[186][88] = 1;
        pixel_data[186][89] = 1;
        pixel_data[186][90] = 1;
        pixel_data[186][91] = 1;
        pixel_data[186][92] = 1;
        pixel_data[186][93] = 1;
        pixel_data[186][94] = 1;
        pixel_data[186][95] = 1;
        pixel_data[186][96] = 1;
        pixel_data[186][97] = 1;
        pixel_data[186][98] = 1;
        pixel_data[186][99] = 1;
        pixel_data[186][100] = 1;
        pixel_data[186][101] = 1;
        pixel_data[186][102] = 1;
        pixel_data[186][103] = 1;
        pixel_data[186][104] = 1;
        pixel_data[186][105] = 1;
        pixel_data[186][106] = 1;
        pixel_data[186][107] = 1;
        pixel_data[186][108] = 1;
        pixel_data[186][109] = 1;
        pixel_data[186][110] = 1;
        pixel_data[186][111] = 1;
        pixel_data[186][112] = 1;
        pixel_data[186][113] = 1;
        pixel_data[186][114] = 1;
        pixel_data[186][115] = 1;
        pixel_data[186][116] = 1;
        pixel_data[186][117] = 1;
        pixel_data[186][118] = 1;
        pixel_data[186][119] = 1;
        pixel_data[186][120] = 1;
        pixel_data[186][121] = 1;
        pixel_data[186][122] = 1;
        pixel_data[186][123] = 1;
        pixel_data[186][124] = 1;
        pixel_data[186][125] = 1;
        pixel_data[186][126] = 1;
        pixel_data[186][127] = 1;
        pixel_data[186][128] = 1;
        pixel_data[186][129] = 1;
        pixel_data[186][130] = 1;
        pixel_data[186][131] = 1;
        pixel_data[186][132] = 1;
        pixel_data[186][133] = 1;
        pixel_data[186][134] = 1;
        pixel_data[186][135] = 1;
        pixel_data[186][136] = 1;
        pixel_data[186][137] = 1;
        pixel_data[186][138] = 1;
        pixel_data[186][139] = 1;
        pixel_data[186][140] = 1;
        pixel_data[186][141] = 1;
        pixel_data[186][142] = 1;
        pixel_data[186][143] = 1;
        pixel_data[186][144] = 1;
        pixel_data[186][145] = 1;
        pixel_data[186][146] = 1;
        pixel_data[186][147] = 1;
        pixel_data[186][148] = 1;
        pixel_data[186][149] = 1;
        pixel_data[186][150] = 1;
        pixel_data[186][151] = 1;
        pixel_data[186][152] = 1;
        pixel_data[186][153] = 1;
        pixel_data[186][154] = 1;
        pixel_data[186][155] = 1;
        pixel_data[186][156] = 1;
        pixel_data[186][157] = 1;
        pixel_data[186][158] = 1;
        pixel_data[186][159] = 1;
        pixel_data[186][160] = 1;
        pixel_data[186][161] = 1;
        pixel_data[186][162] = 1;
        pixel_data[186][163] = 1;
        pixel_data[186][164] = 1;
        pixel_data[186][165] = 1;
        pixel_data[186][166] = 1;
        pixel_data[186][167] = 1;
        pixel_data[186][168] = 1;
        pixel_data[186][169] = 1;
        pixel_data[186][170] = 1;
        pixel_data[186][171] = 1;
        pixel_data[186][172] = 1;
        pixel_data[186][173] = 1;
        pixel_data[186][174] = 1;
        pixel_data[186][175] = 1;
        pixel_data[186][176] = 1;
        pixel_data[186][177] = 1;
        pixel_data[186][178] = 1;
        pixel_data[186][179] = 1;
        pixel_data[186][180] = 1;
        pixel_data[186][181] = 1;
        pixel_data[186][182] = 1;
        pixel_data[186][183] = 1;
        pixel_data[186][184] = 1;
        pixel_data[186][185] = 1;
        pixel_data[186][186] = 1;
        pixel_data[186][187] = 1;
        pixel_data[186][188] = 1;
        pixel_data[186][189] = 5;
        pixel_data[186][190] = 8;
        pixel_data[186][191] = 11;
        pixel_data[186][192] = 11;
        pixel_data[186][193] = 0;
        pixel_data[186][194] = 0;
        pixel_data[186][195] = 0;
        pixel_data[186][196] = 0;
        pixel_data[186][197] = 0;
        pixel_data[186][198] = 0;
        pixel_data[186][199] = 0; // y=186
        pixel_data[187][0] = 0;
        pixel_data[187][1] = 0;
        pixel_data[187][2] = 0;
        pixel_data[187][3] = 10;
        pixel_data[187][4] = 11;
        pixel_data[187][5] = 11;
        pixel_data[187][6] = 7;
        pixel_data[187][7] = 1;
        pixel_data[187][8] = 1;
        pixel_data[187][9] = 1;
        pixel_data[187][10] = 1;
        pixel_data[187][11] = 1;
        pixel_data[187][12] = 1;
        pixel_data[187][13] = 2;
        pixel_data[187][14] = 4;
        pixel_data[187][15] = 4;
        pixel_data[187][16] = 1;
        pixel_data[187][17] = 1;
        pixel_data[187][18] = 1;
        pixel_data[187][19] = 1;
        pixel_data[187][20] = 1;
        pixel_data[187][21] = 1;
        pixel_data[187][22] = 1;
        pixel_data[187][23] = 1;
        pixel_data[187][24] = 1;
        pixel_data[187][25] = 1;
        pixel_data[187][26] = 1;
        pixel_data[187][27] = 1;
        pixel_data[187][28] = 1;
        pixel_data[187][29] = 1;
        pixel_data[187][30] = 1;
        pixel_data[187][31] = 1;
        pixel_data[187][32] = 1;
        pixel_data[187][33] = 1;
        pixel_data[187][34] = 1;
        pixel_data[187][35] = 1;
        pixel_data[187][36] = 1;
        pixel_data[187][37] = 1;
        pixel_data[187][38] = 1;
        pixel_data[187][39] = 1;
        pixel_data[187][40] = 1;
        pixel_data[187][41] = 1;
        pixel_data[187][42] = 1;
        pixel_data[187][43] = 1;
        pixel_data[187][44] = 1;
        pixel_data[187][45] = 1;
        pixel_data[187][46] = 1;
        pixel_data[187][47] = 1;
        pixel_data[187][48] = 1;
        pixel_data[187][49] = 1;
        pixel_data[187][50] = 1;
        pixel_data[187][51] = 1;
        pixel_data[187][52] = 1;
        pixel_data[187][53] = 1;
        pixel_data[187][54] = 1;
        pixel_data[187][55] = 1;
        pixel_data[187][56] = 1;
        pixel_data[187][57] = 1;
        pixel_data[187][58] = 1;
        pixel_data[187][59] = 1;
        pixel_data[187][60] = 1;
        pixel_data[187][61] = 1;
        pixel_data[187][62] = 1;
        pixel_data[187][63] = 1;
        pixel_data[187][64] = 1;
        pixel_data[187][65] = 1;
        pixel_data[187][66] = 1;
        pixel_data[187][67] = 1;
        pixel_data[187][68] = 1;
        pixel_data[187][69] = 1;
        pixel_data[187][70] = 1;
        pixel_data[187][71] = 1;
        pixel_data[187][72] = 1;
        pixel_data[187][73] = 1;
        pixel_data[187][74] = 1;
        pixel_data[187][75] = 1;
        pixel_data[187][76] = 1;
        pixel_data[187][77] = 1;
        pixel_data[187][78] = 1;
        pixel_data[187][79] = 1;
        pixel_data[187][80] = 1;
        pixel_data[187][81] = 1;
        pixel_data[187][82] = 1;
        pixel_data[187][83] = 1;
        pixel_data[187][84] = 1;
        pixel_data[187][85] = 1;
        pixel_data[187][86] = 1;
        pixel_data[187][87] = 1;
        pixel_data[187][88] = 1;
        pixel_data[187][89] = 1;
        pixel_data[187][90] = 1;
        pixel_data[187][91] = 1;
        pixel_data[187][92] = 1;
        pixel_data[187][93] = 1;
        pixel_data[187][94] = 1;
        pixel_data[187][95] = 1;
        pixel_data[187][96] = 1;
        pixel_data[187][97] = 1;
        pixel_data[187][98] = 1;
        pixel_data[187][99] = 1;
        pixel_data[187][100] = 1;
        pixel_data[187][101] = 1;
        pixel_data[187][102] = 1;
        pixel_data[187][103] = 1;
        pixel_data[187][104] = 1;
        pixel_data[187][105] = 1;
        pixel_data[187][106] = 1;
        pixel_data[187][107] = 1;
        pixel_data[187][108] = 1;
        pixel_data[187][109] = 1;
        pixel_data[187][110] = 1;
        pixel_data[187][111] = 1;
        pixel_data[187][112] = 1;
        pixel_data[187][113] = 1;
        pixel_data[187][114] = 1;
        pixel_data[187][115] = 1;
        pixel_data[187][116] = 1;
        pixel_data[187][117] = 1;
        pixel_data[187][118] = 1;
        pixel_data[187][119] = 1;
        pixel_data[187][120] = 1;
        pixel_data[187][121] = 1;
        pixel_data[187][122] = 1;
        pixel_data[187][123] = 1;
        pixel_data[187][124] = 1;
        pixel_data[187][125] = 1;
        pixel_data[187][126] = 1;
        pixel_data[187][127] = 1;
        pixel_data[187][128] = 1;
        pixel_data[187][129] = 1;
        pixel_data[187][130] = 1;
        pixel_data[187][131] = 1;
        pixel_data[187][132] = 1;
        pixel_data[187][133] = 1;
        pixel_data[187][134] = 1;
        pixel_data[187][135] = 1;
        pixel_data[187][136] = 1;
        pixel_data[187][137] = 1;
        pixel_data[187][138] = 1;
        pixel_data[187][139] = 1;
        pixel_data[187][140] = 1;
        pixel_data[187][141] = 1;
        pixel_data[187][142] = 1;
        pixel_data[187][143] = 1;
        pixel_data[187][144] = 1;
        pixel_data[187][145] = 1;
        pixel_data[187][146] = 1;
        pixel_data[187][147] = 1;
        pixel_data[187][148] = 1;
        pixel_data[187][149] = 1;
        pixel_data[187][150] = 1;
        pixel_data[187][151] = 1;
        pixel_data[187][152] = 1;
        pixel_data[187][153] = 1;
        pixel_data[187][154] = 1;
        pixel_data[187][155] = 1;
        pixel_data[187][156] = 1;
        pixel_data[187][157] = 1;
        pixel_data[187][158] = 1;
        pixel_data[187][159] = 1;
        pixel_data[187][160] = 1;
        pixel_data[187][161] = 1;
        pixel_data[187][162] = 1;
        pixel_data[187][163] = 1;
        pixel_data[187][164] = 1;
        pixel_data[187][165] = 1;
        pixel_data[187][166] = 1;
        pixel_data[187][167] = 1;
        pixel_data[187][168] = 1;
        pixel_data[187][169] = 1;
        pixel_data[187][170] = 1;
        pixel_data[187][171] = 1;
        pixel_data[187][172] = 1;
        pixel_data[187][173] = 1;
        pixel_data[187][174] = 1;
        pixel_data[187][175] = 1;
        pixel_data[187][176] = 1;
        pixel_data[187][177] = 1;
        pixel_data[187][178] = 1;
        pixel_data[187][179] = 1;
        pixel_data[187][180] = 1;
        pixel_data[187][181] = 1;
        pixel_data[187][182] = 1;
        pixel_data[187][183] = 1;
        pixel_data[187][184] = 1;
        pixel_data[187][185] = 1;
        pixel_data[187][186] = 1;
        pixel_data[187][187] = 1;
        pixel_data[187][188] = 1;
        pixel_data[187][189] = 4;
        pixel_data[187][190] = 7;
        pixel_data[187][191] = 11;
        pixel_data[187][192] = 11;
        pixel_data[187][193] = 0;
        pixel_data[187][194] = 0;
        pixel_data[187][195] = 0;
        pixel_data[187][196] = 0;
        pixel_data[187][197] = 0;
        pixel_data[187][198] = 0;
        pixel_data[187][199] = 0; // y=187
        pixel_data[188][0] = 0;
        pixel_data[188][1] = 0;
        pixel_data[188][2] = 0;
        pixel_data[188][3] = 0;
        pixel_data[188][4] = 11;
        pixel_data[188][5] = 11;
        pixel_data[188][6] = 8;
        pixel_data[188][7] = 5;
        pixel_data[188][8] = 1;
        pixel_data[188][9] = 1;
        pixel_data[188][10] = 1;
        pixel_data[188][11] = 1;
        pixel_data[188][12] = 1;
        pixel_data[188][13] = 1;
        pixel_data[188][14] = 2;
        pixel_data[188][15] = 4;
        pixel_data[188][16] = 4;
        pixel_data[188][17] = 1;
        pixel_data[188][18] = 1;
        pixel_data[188][19] = 1;
        pixel_data[188][20] = 1;
        pixel_data[188][21] = 1;
        pixel_data[188][22] = 1;
        pixel_data[188][23] = 1;
        pixel_data[188][24] = 1;
        pixel_data[188][25] = 1;
        pixel_data[188][26] = 1;
        pixel_data[188][27] = 1;
        pixel_data[188][28] = 1;
        pixel_data[188][29] = 1;
        pixel_data[188][30] = 1;
        pixel_data[188][31] = 1;
        pixel_data[188][32] = 1;
        pixel_data[188][33] = 1;
        pixel_data[188][34] = 1;
        pixel_data[188][35] = 1;
        pixel_data[188][36] = 1;
        pixel_data[188][37] = 1;
        pixel_data[188][38] = 1;
        pixel_data[188][39] = 1;
        pixel_data[188][40] = 1;
        pixel_data[188][41] = 1;
        pixel_data[188][42] = 1;
        pixel_data[188][43] = 1;
        pixel_data[188][44] = 1;
        pixel_data[188][45] = 1;
        pixel_data[188][46] = 1;
        pixel_data[188][47] = 1;
        pixel_data[188][48] = 1;
        pixel_data[188][49] = 1;
        pixel_data[188][50] = 1;
        pixel_data[188][51] = 1;
        pixel_data[188][52] = 1;
        pixel_data[188][53] = 1;
        pixel_data[188][54] = 1;
        pixel_data[188][55] = 1;
        pixel_data[188][56] = 1;
        pixel_data[188][57] = 1;
        pixel_data[188][58] = 1;
        pixel_data[188][59] = 1;
        pixel_data[188][60] = 1;
        pixel_data[188][61] = 1;
        pixel_data[188][62] = 1;
        pixel_data[188][63] = 1;
        pixel_data[188][64] = 1;
        pixel_data[188][65] = 1;
        pixel_data[188][66] = 1;
        pixel_data[188][67] = 1;
        pixel_data[188][68] = 1;
        pixel_data[188][69] = 1;
        pixel_data[188][70] = 1;
        pixel_data[188][71] = 1;
        pixel_data[188][72] = 1;
        pixel_data[188][73] = 1;
        pixel_data[188][74] = 1;
        pixel_data[188][75] = 1;
        pixel_data[188][76] = 1;
        pixel_data[188][77] = 1;
        pixel_data[188][78] = 1;
        pixel_data[188][79] = 1;
        pixel_data[188][80] = 1;
        pixel_data[188][81] = 1;
        pixel_data[188][82] = 1;
        pixel_data[188][83] = 1;
        pixel_data[188][84] = 1;
        pixel_data[188][85] = 1;
        pixel_data[188][86] = 1;
        pixel_data[188][87] = 1;
        pixel_data[188][88] = 1;
        pixel_data[188][89] = 1;
        pixel_data[188][90] = 1;
        pixel_data[188][91] = 1;
        pixel_data[188][92] = 1;
        pixel_data[188][93] = 1;
        pixel_data[188][94] = 1;
        pixel_data[188][95] = 1;
        pixel_data[188][96] = 1;
        pixel_data[188][97] = 1;
        pixel_data[188][98] = 1;
        pixel_data[188][99] = 1;
        pixel_data[188][100] = 1;
        pixel_data[188][101] = 1;
        pixel_data[188][102] = 1;
        pixel_data[188][103] = 1;
        pixel_data[188][104] = 1;
        pixel_data[188][105] = 1;
        pixel_data[188][106] = 1;
        pixel_data[188][107] = 1;
        pixel_data[188][108] = 1;
        pixel_data[188][109] = 1;
        pixel_data[188][110] = 1;
        pixel_data[188][111] = 1;
        pixel_data[188][112] = 1;
        pixel_data[188][113] = 1;
        pixel_data[188][114] = 1;
        pixel_data[188][115] = 1;
        pixel_data[188][116] = 1;
        pixel_data[188][117] = 1;
        pixel_data[188][118] = 1;
        pixel_data[188][119] = 1;
        pixel_data[188][120] = 1;
        pixel_data[188][121] = 1;
        pixel_data[188][122] = 1;
        pixel_data[188][123] = 1;
        pixel_data[188][124] = 1;
        pixel_data[188][125] = 1;
        pixel_data[188][126] = 1;
        pixel_data[188][127] = 1;
        pixel_data[188][128] = 1;
        pixel_data[188][129] = 1;
        pixel_data[188][130] = 1;
        pixel_data[188][131] = 1;
        pixel_data[188][132] = 1;
        pixel_data[188][133] = 1;
        pixel_data[188][134] = 1;
        pixel_data[188][135] = 1;
        pixel_data[188][136] = 1;
        pixel_data[188][137] = 1;
        pixel_data[188][138] = 1;
        pixel_data[188][139] = 1;
        pixel_data[188][140] = 1;
        pixel_data[188][141] = 1;
        pixel_data[188][142] = 1;
        pixel_data[188][143] = 1;
        pixel_data[188][144] = 1;
        pixel_data[188][145] = 1;
        pixel_data[188][146] = 1;
        pixel_data[188][147] = 1;
        pixel_data[188][148] = 1;
        pixel_data[188][149] = 1;
        pixel_data[188][150] = 1;
        pixel_data[188][151] = 1;
        pixel_data[188][152] = 1;
        pixel_data[188][153] = 1;
        pixel_data[188][154] = 1;
        pixel_data[188][155] = 1;
        pixel_data[188][156] = 1;
        pixel_data[188][157] = 1;
        pixel_data[188][158] = 1;
        pixel_data[188][159] = 1;
        pixel_data[188][160] = 1;
        pixel_data[188][161] = 1;
        pixel_data[188][162] = 1;
        pixel_data[188][163] = 1;
        pixel_data[188][164] = 1;
        pixel_data[188][165] = 1;
        pixel_data[188][166] = 1;
        pixel_data[188][167] = 1;
        pixel_data[188][168] = 1;
        pixel_data[188][169] = 1;
        pixel_data[188][170] = 1;
        pixel_data[188][171] = 1;
        pixel_data[188][172] = 1;
        pixel_data[188][173] = 1;
        pixel_data[188][174] = 1;
        pixel_data[188][175] = 1;
        pixel_data[188][176] = 1;
        pixel_data[188][177] = 1;
        pixel_data[188][178] = 1;
        pixel_data[188][179] = 1;
        pixel_data[188][180] = 1;
        pixel_data[188][181] = 1;
        pixel_data[188][182] = 1;
        pixel_data[188][183] = 1;
        pixel_data[188][184] = 1;
        pixel_data[188][185] = 1;
        pixel_data[188][186] = 1;
        pixel_data[188][187] = 1;
        pixel_data[188][188] = 1;
        pixel_data[188][189] = 5;
        pixel_data[188][190] = 8;
        pixel_data[188][191] = 11;
        pixel_data[188][192] = 11;
        pixel_data[188][193] = 0;
        pixel_data[188][194] = 0;
        pixel_data[188][195] = 0;
        pixel_data[188][196] = 0;
        pixel_data[188][197] = 0;
        pixel_data[188][198] = 0;
        pixel_data[188][199] = 0; // y=188
        pixel_data[189][0] = 0;
        pixel_data[189][1] = 0;
        pixel_data[189][2] = 0;
        pixel_data[189][3] = 0;
        pixel_data[189][4] = 11;
        pixel_data[189][5] = 11;
        pixel_data[189][6] = 9;
        pixel_data[189][7] = 7;
        pixel_data[189][8] = 1;
        pixel_data[189][9] = 1;
        pixel_data[189][10] = 1;
        pixel_data[189][11] = 1;
        pixel_data[189][12] = 1;
        pixel_data[189][13] = 1;
        pixel_data[189][14] = 1;
        pixel_data[189][15] = 4;
        pixel_data[189][16] = 4;
        pixel_data[189][17] = 2;
        pixel_data[189][18] = 1;
        pixel_data[189][19] = 1;
        pixel_data[189][20] = 1;
        pixel_data[189][21] = 1;
        pixel_data[189][22] = 1;
        pixel_data[189][23] = 1;
        pixel_data[189][24] = 1;
        pixel_data[189][25] = 1;
        pixel_data[189][26] = 1;
        pixel_data[189][27] = 1;
        pixel_data[189][28] = 1;
        pixel_data[189][29] = 1;
        pixel_data[189][30] = 1;
        pixel_data[189][31] = 1;
        pixel_data[189][32] = 1;
        pixel_data[189][33] = 1;
        pixel_data[189][34] = 1;
        pixel_data[189][35] = 1;
        pixel_data[189][36] = 1;
        pixel_data[189][37] = 1;
        pixel_data[189][38] = 1;
        pixel_data[189][39] = 1;
        pixel_data[189][40] = 1;
        pixel_data[189][41] = 1;
        pixel_data[189][42] = 1;
        pixel_data[189][43] = 1;
        pixel_data[189][44] = 1;
        pixel_data[189][45] = 1;
        pixel_data[189][46] = 1;
        pixel_data[189][47] = 1;
        pixel_data[189][48] = 1;
        pixel_data[189][49] = 1;
        pixel_data[189][50] = 1;
        pixel_data[189][51] = 1;
        pixel_data[189][52] = 1;
        pixel_data[189][53] = 1;
        pixel_data[189][54] = 1;
        pixel_data[189][55] = 1;
        pixel_data[189][56] = 1;
        pixel_data[189][57] = 1;
        pixel_data[189][58] = 1;
        pixel_data[189][59] = 1;
        pixel_data[189][60] = 1;
        pixel_data[189][61] = 1;
        pixel_data[189][62] = 1;
        pixel_data[189][63] = 1;
        pixel_data[189][64] = 1;
        pixel_data[189][65] = 1;
        pixel_data[189][66] = 1;
        pixel_data[189][67] = 1;
        pixel_data[189][68] = 1;
        pixel_data[189][69] = 1;
        pixel_data[189][70] = 1;
        pixel_data[189][71] = 1;
        pixel_data[189][72] = 1;
        pixel_data[189][73] = 1;
        pixel_data[189][74] = 1;
        pixel_data[189][75] = 1;
        pixel_data[189][76] = 1;
        pixel_data[189][77] = 1;
        pixel_data[189][78] = 1;
        pixel_data[189][79] = 1;
        pixel_data[189][80] = 1;
        pixel_data[189][81] = 1;
        pixel_data[189][82] = 1;
        pixel_data[189][83] = 1;
        pixel_data[189][84] = 1;
        pixel_data[189][85] = 1;
        pixel_data[189][86] = 1;
        pixel_data[189][87] = 1;
        pixel_data[189][88] = 1;
        pixel_data[189][89] = 1;
        pixel_data[189][90] = 1;
        pixel_data[189][91] = 1;
        pixel_data[189][92] = 1;
        pixel_data[189][93] = 1;
        pixel_data[189][94] = 1;
        pixel_data[189][95] = 1;
        pixel_data[189][96] = 1;
        pixel_data[189][97] = 1;
        pixel_data[189][98] = 1;
        pixel_data[189][99] = 1;
        pixel_data[189][100] = 1;
        pixel_data[189][101] = 1;
        pixel_data[189][102] = 1;
        pixel_data[189][103] = 1;
        pixel_data[189][104] = 1;
        pixel_data[189][105] = 1;
        pixel_data[189][106] = 1;
        pixel_data[189][107] = 1;
        pixel_data[189][108] = 1;
        pixel_data[189][109] = 1;
        pixel_data[189][110] = 1;
        pixel_data[189][111] = 1;
        pixel_data[189][112] = 1;
        pixel_data[189][113] = 1;
        pixel_data[189][114] = 1;
        pixel_data[189][115] = 1;
        pixel_data[189][116] = 1;
        pixel_data[189][117] = 1;
        pixel_data[189][118] = 1;
        pixel_data[189][119] = 1;
        pixel_data[189][120] = 1;
        pixel_data[189][121] = 1;
        pixel_data[189][122] = 1;
        pixel_data[189][123] = 1;
        pixel_data[189][124] = 1;
        pixel_data[189][125] = 1;
        pixel_data[189][126] = 1;
        pixel_data[189][127] = 1;
        pixel_data[189][128] = 1;
        pixel_data[189][129] = 1;
        pixel_data[189][130] = 1;
        pixel_data[189][131] = 1;
        pixel_data[189][132] = 1;
        pixel_data[189][133] = 1;
        pixel_data[189][134] = 1;
        pixel_data[189][135] = 1;
        pixel_data[189][136] = 1;
        pixel_data[189][137] = 1;
        pixel_data[189][138] = 1;
        pixel_data[189][139] = 1;
        pixel_data[189][140] = 1;
        pixel_data[189][141] = 1;
        pixel_data[189][142] = 1;
        pixel_data[189][143] = 1;
        pixel_data[189][144] = 1;
        pixel_data[189][145] = 1;
        pixel_data[189][146] = 1;
        pixel_data[189][147] = 1;
        pixel_data[189][148] = 1;
        pixel_data[189][149] = 1;
        pixel_data[189][150] = 1;
        pixel_data[189][151] = 1;
        pixel_data[189][152] = 1;
        pixel_data[189][153] = 1;
        pixel_data[189][154] = 1;
        pixel_data[189][155] = 1;
        pixel_data[189][156] = 1;
        pixel_data[189][157] = 1;
        pixel_data[189][158] = 1;
        pixel_data[189][159] = 1;
        pixel_data[189][160] = 1;
        pixel_data[189][161] = 1;
        pixel_data[189][162] = 1;
        pixel_data[189][163] = 1;
        pixel_data[189][164] = 1;
        pixel_data[189][165] = 1;
        pixel_data[189][166] = 1;
        pixel_data[189][167] = 1;
        pixel_data[189][168] = 1;
        pixel_data[189][169] = 1;
        pixel_data[189][170] = 1;
        pixel_data[189][171] = 1;
        pixel_data[189][172] = 1;
        pixel_data[189][173] = 1;
        pixel_data[189][174] = 1;
        pixel_data[189][175] = 1;
        pixel_data[189][176] = 1;
        pixel_data[189][177] = 1;
        pixel_data[189][178] = 1;
        pixel_data[189][179] = 1;
        pixel_data[189][180] = 1;
        pixel_data[189][181] = 1;
        pixel_data[189][182] = 1;
        pixel_data[189][183] = 1;
        pixel_data[189][184] = 1;
        pixel_data[189][185] = 1;
        pixel_data[189][186] = 1;
        pixel_data[189][187] = 1;
        pixel_data[189][188] = 1;
        pixel_data[189][189] = 7;
        pixel_data[189][190] = 9;
        pixel_data[189][191] = 11;
        pixel_data[189][192] = 11;
        pixel_data[189][193] = 0;
        pixel_data[189][194] = 0;
        pixel_data[189][195] = 0;
        pixel_data[189][196] = 0;
        pixel_data[189][197] = 0;
        pixel_data[189][198] = 0;
        pixel_data[189][199] = 0; // y=189
        pixel_data[190][0] = 0;
        pixel_data[190][1] = 0;
        pixel_data[190][2] = 0;
        pixel_data[190][3] = 0;
        pixel_data[190][4] = 0;
        pixel_data[190][5] = 11;
        pixel_data[190][6] = 11;
        pixel_data[190][7] = 8;
        pixel_data[190][8] = 6;
        pixel_data[190][9] = 1;
        pixel_data[190][10] = 1;
        pixel_data[190][11] = 1;
        pixel_data[190][12] = 1;
        pixel_data[190][13] = 1;
        pixel_data[190][14] = 1;
        pixel_data[190][15] = 4;
        pixel_data[190][16] = 4;
        pixel_data[190][17] = 4;
        pixel_data[190][18] = 1;
        pixel_data[190][19] = 1;
        pixel_data[190][20] = 1;
        pixel_data[190][21] = 1;
        pixel_data[190][22] = 1;
        pixel_data[190][23] = 1;
        pixel_data[190][24] = 1;
        pixel_data[190][25] = 1;
        pixel_data[190][26] = 1;
        pixel_data[190][27] = 1;
        pixel_data[190][28] = 1;
        pixel_data[190][29] = 1;
        pixel_data[190][30] = 1;
        pixel_data[190][31] = 1;
        pixel_data[190][32] = 1;
        pixel_data[190][33] = 1;
        pixel_data[190][34] = 1;
        pixel_data[190][35] = 1;
        pixel_data[190][36] = 1;
        pixel_data[190][37] = 4;
        pixel_data[190][38] = 4;
        pixel_data[190][39] = 2;
        pixel_data[190][40] = 1;
        pixel_data[190][41] = 1;
        pixel_data[190][42] = 1;
        pixel_data[190][43] = 1;
        pixel_data[190][44] = 1;
        pixel_data[190][45] = 1;
        pixel_data[190][46] = 1;
        pixel_data[190][47] = 1;
        pixel_data[190][48] = 1;
        pixel_data[190][49] = 1;
        pixel_data[190][50] = 1;
        pixel_data[190][51] = 1;
        pixel_data[190][52] = 1;
        pixel_data[190][53] = 1;
        pixel_data[190][54] = 1;
        pixel_data[190][55] = 1;
        pixel_data[190][56] = 1;
        pixel_data[190][57] = 1;
        pixel_data[190][58] = 1;
        pixel_data[190][59] = 1;
        pixel_data[190][60] = 1;
        pixel_data[190][61] = 1;
        pixel_data[190][62] = 1;
        pixel_data[190][63] = 1;
        pixel_data[190][64] = 1;
        pixel_data[190][65] = 1;
        pixel_data[190][66] = 1;
        pixel_data[190][67] = 1;
        pixel_data[190][68] = 1;
        pixel_data[190][69] = 1;
        pixel_data[190][70] = 1;
        pixel_data[190][71] = 1;
        pixel_data[190][72] = 1;
        pixel_data[190][73] = 1;
        pixel_data[190][74] = 1;
        pixel_data[190][75] = 1;
        pixel_data[190][76] = 1;
        pixel_data[190][77] = 1;
        pixel_data[190][78] = 1;
        pixel_data[190][79] = 1;
        pixel_data[190][80] = 1;
        pixel_data[190][81] = 1;
        pixel_data[190][82] = 1;
        pixel_data[190][83] = 1;
        pixel_data[190][84] = 1;
        pixel_data[190][85] = 1;
        pixel_data[190][86] = 1;
        pixel_data[190][87] = 1;
        pixel_data[190][88] = 1;
        pixel_data[190][89] = 1;
        pixel_data[190][90] = 1;
        pixel_data[190][91] = 1;
        pixel_data[190][92] = 1;
        pixel_data[190][93] = 1;
        pixel_data[190][94] = 1;
        pixel_data[190][95] = 1;
        pixel_data[190][96] = 1;
        pixel_data[190][97] = 1;
        pixel_data[190][98] = 1;
        pixel_data[190][99] = 1;
        pixel_data[190][100] = 1;
        pixel_data[190][101] = 1;
        pixel_data[190][102] = 1;
        pixel_data[190][103] = 1;
        pixel_data[190][104] = 1;
        pixel_data[190][105] = 1;
        pixel_data[190][106] = 1;
        pixel_data[190][107] = 1;
        pixel_data[190][108] = 1;
        pixel_data[190][109] = 1;
        pixel_data[190][110] = 1;
        pixel_data[190][111] = 1;
        pixel_data[190][112] = 1;
        pixel_data[190][113] = 1;
        pixel_data[190][114] = 1;
        pixel_data[190][115] = 1;
        pixel_data[190][116] = 1;
        pixel_data[190][117] = 1;
        pixel_data[190][118] = 1;
        pixel_data[190][119] = 1;
        pixel_data[190][120] = 1;
        pixel_data[190][121] = 1;
        pixel_data[190][122] = 1;
        pixel_data[190][123] = 1;
        pixel_data[190][124] = 1;
        pixel_data[190][125] = 1;
        pixel_data[190][126] = 1;
        pixel_data[190][127] = 1;
        pixel_data[190][128] = 1;
        pixel_data[190][129] = 1;
        pixel_data[190][130] = 1;
        pixel_data[190][131] = 1;
        pixel_data[190][132] = 1;
        pixel_data[190][133] = 1;
        pixel_data[190][134] = 1;
        pixel_data[190][135] = 1;
        pixel_data[190][136] = 1;
        pixel_data[190][137] = 1;
        pixel_data[190][138] = 1;
        pixel_data[190][139] = 1;
        pixel_data[190][140] = 1;
        pixel_data[190][141] = 1;
        pixel_data[190][142] = 1;
        pixel_data[190][143] = 1;
        pixel_data[190][144] = 1;
        pixel_data[190][145] = 1;
        pixel_data[190][146] = 1;
        pixel_data[190][147] = 1;
        pixel_data[190][148] = 1;
        pixel_data[190][149] = 1;
        pixel_data[190][150] = 1;
        pixel_data[190][151] = 1;
        pixel_data[190][152] = 1;
        pixel_data[190][153] = 1;
        pixel_data[190][154] = 1;
        pixel_data[190][155] = 1;
        pixel_data[190][156] = 1;
        pixel_data[190][157] = 1;
        pixel_data[190][158] = 1;
        pixel_data[190][159] = 1;
        pixel_data[190][160] = 1;
        pixel_data[190][161] = 1;
        pixel_data[190][162] = 1;
        pixel_data[190][163] = 1;
        pixel_data[190][164] = 1;
        pixel_data[190][165] = 1;
        pixel_data[190][166] = 1;
        pixel_data[190][167] = 1;
        pixel_data[190][168] = 1;
        pixel_data[190][169] = 1;
        pixel_data[190][170] = 1;
        pixel_data[190][171] = 1;
        pixel_data[190][172] = 1;
        pixel_data[190][173] = 1;
        pixel_data[190][174] = 1;
        pixel_data[190][175] = 1;
        pixel_data[190][176] = 1;
        pixel_data[190][177] = 1;
        pixel_data[190][178] = 1;
        pixel_data[190][179] = 1;
        pixel_data[190][180] = 1;
        pixel_data[190][181] = 1;
        pixel_data[190][182] = 1;
        pixel_data[190][183] = 1;
        pixel_data[190][184] = 1;
        pixel_data[190][185] = 1;
        pixel_data[190][186] = 1;
        pixel_data[190][187] = 1;
        pixel_data[190][188] = 6;
        pixel_data[190][189] = 8;
        pixel_data[190][190] = 11;
        pixel_data[190][191] = 11;
        pixel_data[190][192] = 0;
        pixel_data[190][193] = 0;
        pixel_data[190][194] = 0;
        pixel_data[190][195] = 0;
        pixel_data[190][196] = 0;
        pixel_data[190][197] = 0;
        pixel_data[190][198] = 0;
        pixel_data[190][199] = 0; // y=190
        pixel_data[191][0] = 0;
        pixel_data[191][1] = 0;
        pixel_data[191][2] = 0;
        pixel_data[191][3] = 0;
        pixel_data[191][4] = 0;
        pixel_data[191][5] = 0;
        pixel_data[191][6] = 11;
        pixel_data[191][7] = 11;
        pixel_data[191][8] = 8;
        pixel_data[191][9] = 5;
        pixel_data[191][10] = 1;
        pixel_data[191][11] = 1;
        pixel_data[191][12] = 1;
        pixel_data[191][13] = 1;
        pixel_data[191][14] = 1;
        pixel_data[191][15] = 1;
        pixel_data[191][16] = 4;
        pixel_data[191][17] = 4;
        pixel_data[191][18] = 2;
        pixel_data[191][19] = 1;
        pixel_data[191][20] = 1;
        pixel_data[191][21] = 1;
        pixel_data[191][22] = 1;
        pixel_data[191][23] = 1;
        pixel_data[191][24] = 1;
        pixel_data[191][25] = 1;
        pixel_data[191][26] = 1;
        pixel_data[191][27] = 1;
        pixel_data[191][28] = 1;
        pixel_data[191][29] = 1;
        pixel_data[191][30] = 1;
        pixel_data[191][31] = 1;
        pixel_data[191][32] = 1;
        pixel_data[191][33] = 1;
        pixel_data[191][34] = 1;
        pixel_data[191][35] = 1;
        pixel_data[191][36] = 4;
        pixel_data[191][37] = 4;
        pixel_data[191][38] = 2;
        pixel_data[191][39] = 1;
        pixel_data[191][40] = 1;
        pixel_data[191][41] = 1;
        pixel_data[191][42] = 1;
        pixel_data[191][43] = 1;
        pixel_data[191][44] = 1;
        pixel_data[191][45] = 1;
        pixel_data[191][46] = 1;
        pixel_data[191][47] = 1;
        pixel_data[191][48] = 1;
        pixel_data[191][49] = 1;
        pixel_data[191][50] = 1;
        pixel_data[191][51] = 1;
        pixel_data[191][52] = 1;
        pixel_data[191][53] = 1;
        pixel_data[191][54] = 1;
        pixel_data[191][55] = 1;
        pixel_data[191][56] = 1;
        pixel_data[191][57] = 1;
        pixel_data[191][58] = 1;
        pixel_data[191][59] = 1;
        pixel_data[191][60] = 1;
        pixel_data[191][61] = 1;
        pixel_data[191][62] = 1;
        pixel_data[191][63] = 1;
        pixel_data[191][64] = 1;
        pixel_data[191][65] = 1;
        pixel_data[191][66] = 1;
        pixel_data[191][67] = 1;
        pixel_data[191][68] = 1;
        pixel_data[191][69] = 1;
        pixel_data[191][70] = 1;
        pixel_data[191][71] = 1;
        pixel_data[191][72] = 1;
        pixel_data[191][73] = 1;
        pixel_data[191][74] = 1;
        pixel_data[191][75] = 1;
        pixel_data[191][76] = 1;
        pixel_data[191][77] = 1;
        pixel_data[191][78] = 1;
        pixel_data[191][79] = 1;
        pixel_data[191][80] = 1;
        pixel_data[191][81] = 1;
        pixel_data[191][82] = 1;
        pixel_data[191][83] = 1;
        pixel_data[191][84] = 1;
        pixel_data[191][85] = 1;
        pixel_data[191][86] = 1;
        pixel_data[191][87] = 1;
        pixel_data[191][88] = 1;
        pixel_data[191][89] = 1;
        pixel_data[191][90] = 1;
        pixel_data[191][91] = 1;
        pixel_data[191][92] = 1;
        pixel_data[191][93] = 1;
        pixel_data[191][94] = 1;
        pixel_data[191][95] = 1;
        pixel_data[191][96] = 1;
        pixel_data[191][97] = 1;
        pixel_data[191][98] = 1;
        pixel_data[191][99] = 1;
        pixel_data[191][100] = 1;
        pixel_data[191][101] = 1;
        pixel_data[191][102] = 1;
        pixel_data[191][103] = 1;
        pixel_data[191][104] = 1;
        pixel_data[191][105] = 1;
        pixel_data[191][106] = 1;
        pixel_data[191][107] = 1;
        pixel_data[191][108] = 1;
        pixel_data[191][109] = 1;
        pixel_data[191][110] = 1;
        pixel_data[191][111] = 1;
        pixel_data[191][112] = 1;
        pixel_data[191][113] = 1;
        pixel_data[191][114] = 1;
        pixel_data[191][115] = 1;
        pixel_data[191][116] = 1;
        pixel_data[191][117] = 1;
        pixel_data[191][118] = 1;
        pixel_data[191][119] = 1;
        pixel_data[191][120] = 1;
        pixel_data[191][121] = 1;
        pixel_data[191][122] = 1;
        pixel_data[191][123] = 1;
        pixel_data[191][124] = 1;
        pixel_data[191][125] = 1;
        pixel_data[191][126] = 1;
        pixel_data[191][127] = 1;
        pixel_data[191][128] = 1;
        pixel_data[191][129] = 1;
        pixel_data[191][130] = 1;
        pixel_data[191][131] = 1;
        pixel_data[191][132] = 1;
        pixel_data[191][133] = 1;
        pixel_data[191][134] = 1;
        pixel_data[191][135] = 1;
        pixel_data[191][136] = 1;
        pixel_data[191][137] = 1;
        pixel_data[191][138] = 1;
        pixel_data[191][139] = 1;
        pixel_data[191][140] = 1;
        pixel_data[191][141] = 1;
        pixel_data[191][142] = 1;
        pixel_data[191][143] = 1;
        pixel_data[191][144] = 1;
        pixel_data[191][145] = 1;
        pixel_data[191][146] = 1;
        pixel_data[191][147] = 1;
        pixel_data[191][148] = 1;
        pixel_data[191][149] = 1;
        pixel_data[191][150] = 1;
        pixel_data[191][151] = 1;
        pixel_data[191][152] = 1;
        pixel_data[191][153] = 1;
        pixel_data[191][154] = 1;
        pixel_data[191][155] = 1;
        pixel_data[191][156] = 1;
        pixel_data[191][157] = 1;
        pixel_data[191][158] = 1;
        pixel_data[191][159] = 1;
        pixel_data[191][160] = 1;
        pixel_data[191][161] = 1;
        pixel_data[191][162] = 1;
        pixel_data[191][163] = 1;
        pixel_data[191][164] = 1;
        pixel_data[191][165] = 1;
        pixel_data[191][166] = 1;
        pixel_data[191][167] = 1;
        pixel_data[191][168] = 1;
        pixel_data[191][169] = 1;
        pixel_data[191][170] = 1;
        pixel_data[191][171] = 1;
        pixel_data[191][172] = 1;
        pixel_data[191][173] = 1;
        pixel_data[191][174] = 1;
        pixel_data[191][175] = 1;
        pixel_data[191][176] = 1;
        pixel_data[191][177] = 1;
        pixel_data[191][178] = 1;
        pixel_data[191][179] = 1;
        pixel_data[191][180] = 1;
        pixel_data[191][181] = 1;
        pixel_data[191][182] = 1;
        pixel_data[191][183] = 1;
        pixel_data[191][184] = 1;
        pixel_data[191][185] = 5;
        pixel_data[191][186] = 8;
        pixel_data[191][187] = 11;
        pixel_data[191][188] = 11;
        pixel_data[191][189] = 11;
        pixel_data[191][190] = 11;
        pixel_data[191][191] = 0;
        pixel_data[191][192] = 0;
        pixel_data[191][193] = 0;
        pixel_data[191][194] = 0;
        pixel_data[191][195] = 0;
        pixel_data[191][196] = 0;
        pixel_data[191][197] = 0;
        pixel_data[191][198] = 0;
        pixel_data[191][199] = 0; // y=191
        pixel_data[192][0] = 0;
        pixel_data[192][1] = 0;
        pixel_data[192][2] = 0;
        pixel_data[192][3] = 0;
        pixel_data[192][4] = 0;
        pixel_data[192][5] = 0;
        pixel_data[192][6] = 10;
        pixel_data[192][7] = 11;
        pixel_data[192][8] = 9;
        pixel_data[192][9] = 7;
        pixel_data[192][10] = 1;
        pixel_data[192][11] = 1;
        pixel_data[192][12] = 1;
        pixel_data[192][13] = 1;
        pixel_data[192][14] = 1;
        pixel_data[192][15] = 1;
        pixel_data[192][16] = 2;
        pixel_data[192][17] = 4;
        pixel_data[192][18] = 4;
        pixel_data[192][19] = 1;
        pixel_data[192][20] = 1;
        pixel_data[192][21] = 1;
        pixel_data[192][22] = 1;
        pixel_data[192][23] = 1;
        pixel_data[192][24] = 1;
        pixel_data[192][25] = 1;
        pixel_data[192][26] = 1;
        pixel_data[192][27] = 1;
        pixel_data[192][28] = 1;
        pixel_data[192][29] = 1;
        pixel_data[192][30] = 1;
        pixel_data[192][31] = 1;
        pixel_data[192][32] = 1;
        pixel_data[192][33] = 1;
        pixel_data[192][34] = 1;
        pixel_data[192][35] = 1;
        pixel_data[192][36] = 4;
        pixel_data[192][37] = 4;
        pixel_data[192][38] = 2;
        pixel_data[192][39] = 1;
        pixel_data[192][40] = 1;
        pixel_data[192][41] = 1;
        pixel_data[192][42] = 1;
        pixel_data[192][43] = 1;
        pixel_data[192][44] = 5;
        pixel_data[192][45] = 7;
        pixel_data[192][46] = 8;
        pixel_data[192][47] = 5;
        pixel_data[192][48] = 1;
        pixel_data[192][49] = 1;
        pixel_data[192][50] = 1;
        pixel_data[192][51] = 1;
        pixel_data[192][52] = 1;
        pixel_data[192][53] = 1;
        pixel_data[192][54] = 1;
        pixel_data[192][55] = 1;
        pixel_data[192][56] = 1;
        pixel_data[192][57] = 1;
        pixel_data[192][58] = 1;
        pixel_data[192][59] = 1;
        pixel_data[192][60] = 1;
        pixel_data[192][61] = 1;
        pixel_data[192][62] = 1;
        pixel_data[192][63] = 1;
        pixel_data[192][64] = 1;
        pixel_data[192][65] = 1;
        pixel_data[192][66] = 1;
        pixel_data[192][67] = 1;
        pixel_data[192][68] = 1;
        pixel_data[192][69] = 1;
        pixel_data[192][70] = 1;
        pixel_data[192][71] = 1;
        pixel_data[192][72] = 1;
        pixel_data[192][73] = 1;
        pixel_data[192][74] = 1;
        pixel_data[192][75] = 1;
        pixel_data[192][76] = 1;
        pixel_data[192][77] = 1;
        pixel_data[192][78] = 1;
        pixel_data[192][79] = 1;
        pixel_data[192][80] = 1;
        pixel_data[192][81] = 1;
        pixel_data[192][82] = 1;
        pixel_data[192][83] = 1;
        pixel_data[192][84] = 1;
        pixel_data[192][85] = 1;
        pixel_data[192][86] = 1;
        pixel_data[192][87] = 1;
        pixel_data[192][88] = 1;
        pixel_data[192][89] = 1;
        pixel_data[192][90] = 1;
        pixel_data[192][91] = 1;
        pixel_data[192][92] = 1;
        pixel_data[192][93] = 1;
        pixel_data[192][94] = 1;
        pixel_data[192][95] = 1;
        pixel_data[192][96] = 1;
        pixel_data[192][97] = 1;
        pixel_data[192][98] = 1;
        pixel_data[192][99] = 1;
        pixel_data[192][100] = 1;
        pixel_data[192][101] = 1;
        pixel_data[192][102] = 1;
        pixel_data[192][103] = 1;
        pixel_data[192][104] = 1;
        pixel_data[192][105] = 1;
        pixel_data[192][106] = 1;
        pixel_data[192][107] = 1;
        pixel_data[192][108] = 1;
        pixel_data[192][109] = 1;
        pixel_data[192][110] = 1;
        pixel_data[192][111] = 1;
        pixel_data[192][112] = 1;
        pixel_data[192][113] = 1;
        pixel_data[192][114] = 1;
        pixel_data[192][115] = 1;
        pixel_data[192][116] = 1;
        pixel_data[192][117] = 1;
        pixel_data[192][118] = 1;
        pixel_data[192][119] = 1;
        pixel_data[192][120] = 1;
        pixel_data[192][121] = 1;
        pixel_data[192][122] = 1;
        pixel_data[192][123] = 1;
        pixel_data[192][124] = 1;
        pixel_data[192][125] = 1;
        pixel_data[192][126] = 1;
        pixel_data[192][127] = 1;
        pixel_data[192][128] = 1;
        pixel_data[192][129] = 1;
        pixel_data[192][130] = 1;
        pixel_data[192][131] = 1;
        pixel_data[192][132] = 1;
        pixel_data[192][133] = 1;
        pixel_data[192][134] = 1;
        pixel_data[192][135] = 1;
        pixel_data[192][136] = 1;
        pixel_data[192][137] = 1;
        pixel_data[192][138] = 1;
        pixel_data[192][139] = 1;
        pixel_data[192][140] = 1;
        pixel_data[192][141] = 1;
        pixel_data[192][142] = 1;
        pixel_data[192][143] = 1;
        pixel_data[192][144] = 1;
        pixel_data[192][145] = 1;
        pixel_data[192][146] = 1;
        pixel_data[192][147] = 1;
        pixel_data[192][148] = 1;
        pixel_data[192][149] = 1;
        pixel_data[192][150] = 1;
        pixel_data[192][151] = 1;
        pixel_data[192][152] = 1;
        pixel_data[192][153] = 1;
        pixel_data[192][154] = 1;
        pixel_data[192][155] = 1;
        pixel_data[192][156] = 1;
        pixel_data[192][157] = 1;
        pixel_data[192][158] = 1;
        pixel_data[192][159] = 1;
        pixel_data[192][160] = 1;
        pixel_data[192][161] = 1;
        pixel_data[192][162] = 1;
        pixel_data[192][163] = 1;
        pixel_data[192][164] = 1;
        pixel_data[192][165] = 1;
        pixel_data[192][166] = 1;
        pixel_data[192][167] = 1;
        pixel_data[192][168] = 1;
        pixel_data[192][169] = 1;
        pixel_data[192][170] = 1;
        pixel_data[192][171] = 1;
        pixel_data[192][172] = 1;
        pixel_data[192][173] = 1;
        pixel_data[192][174] = 1;
        pixel_data[192][175] = 1;
        pixel_data[192][176] = 1;
        pixel_data[192][177] = 1;
        pixel_data[192][178] = 1;
        pixel_data[192][179] = 1;
        pixel_data[192][180] = 1;
        pixel_data[192][181] = 1;
        pixel_data[192][182] = 1;
        pixel_data[192][183] = 5;
        pixel_data[192][184] = 8;
        pixel_data[192][185] = 9;
        pixel_data[192][186] = 11;
        pixel_data[192][187] = 11;
        pixel_data[192][188] = 0;
        pixel_data[192][189] = 0;
        pixel_data[192][190] = 0;
        pixel_data[192][191] = 0;
        pixel_data[192][192] = 0;
        pixel_data[192][193] = 0;
        pixel_data[192][194] = 0;
        pixel_data[192][195] = 0;
        pixel_data[192][196] = 0;
        pixel_data[192][197] = 0;
        pixel_data[192][198] = 0;
        pixel_data[192][199] = 0; // y=192
        pixel_data[193][0] = 0;
        pixel_data[193][1] = 0;
        pixel_data[193][2] = 0;
        pixel_data[193][3] = 0;
        pixel_data[193][4] = 0;
        pixel_data[193][5] = 0;
        pixel_data[193][6] = 0;
        pixel_data[193][7] = 11;
        pixel_data[193][8] = 11;
        pixel_data[193][9] = 9;
        pixel_data[193][10] = 6;
        pixel_data[193][11] = 1;
        pixel_data[193][12] = 1;
        pixel_data[193][13] = 1;
        pixel_data[193][14] = 1;
        pixel_data[193][15] = 1;
        pixel_data[193][16] = 1;
        pixel_data[193][17] = 4;
        pixel_data[193][18] = 4;
        pixel_data[193][19] = 4;
        pixel_data[193][20] = 1;
        pixel_data[193][21] = 1;
        pixel_data[193][22] = 1;
        pixel_data[193][23] = 1;
        pixel_data[193][24] = 1;
        pixel_data[193][25] = 1;
        pixel_data[193][26] = 1;
        pixel_data[193][27] = 1;
        pixel_data[193][28] = 1;
        pixel_data[193][29] = 1;
        pixel_data[193][30] = 1;
        pixel_data[193][31] = 1;
        pixel_data[193][32] = 1;
        pixel_data[193][33] = 1;
        pixel_data[193][34] = 1;
        pixel_data[193][35] = 1;
        pixel_data[193][36] = 4;
        pixel_data[193][37] = 4;
        pixel_data[193][38] = 2;
        pixel_data[193][39] = 1;
        pixel_data[193][40] = 1;
        pixel_data[193][41] = 1;
        pixel_data[193][42] = 5;
        pixel_data[193][43] = 7;
        pixel_data[193][44] = 9;
        pixel_data[193][45] = 11;
        pixel_data[193][46] = 11;
        pixel_data[193][47] = 8;
        pixel_data[193][48] = 5;
        pixel_data[193][49] = 1;
        pixel_data[193][50] = 1;
        pixel_data[193][51] = 1;
        pixel_data[193][52] = 1;
        pixel_data[193][53] = 1;
        pixel_data[193][54] = 1;
        pixel_data[193][55] = 1;
        pixel_data[193][56] = 1;
        pixel_data[193][57] = 1;
        pixel_data[193][58] = 1;
        pixel_data[193][59] = 1;
        pixel_data[193][60] = 1;
        pixel_data[193][61] = 1;
        pixel_data[193][62] = 1;
        pixel_data[193][63] = 1;
        pixel_data[193][64] = 1;
        pixel_data[193][65] = 1;
        pixel_data[193][66] = 1;
        pixel_data[193][67] = 1;
        pixel_data[193][68] = 1;
        pixel_data[193][69] = 1;
        pixel_data[193][70] = 1;
        pixel_data[193][71] = 1;
        pixel_data[193][72] = 1;
        pixel_data[193][73] = 1;
        pixel_data[193][74] = 1;
        pixel_data[193][75] = 1;
        pixel_data[193][76] = 1;
        pixel_data[193][77] = 1;
        pixel_data[193][78] = 1;
        pixel_data[193][79] = 1;
        pixel_data[193][80] = 1;
        pixel_data[193][81] = 1;
        pixel_data[193][82] = 1;
        pixel_data[193][83] = 1;
        pixel_data[193][84] = 1;
        pixel_data[193][85] = 1;
        pixel_data[193][86] = 1;
        pixel_data[193][87] = 1;
        pixel_data[193][88] = 1;
        pixel_data[193][89] = 1;
        pixel_data[193][90] = 1;
        pixel_data[193][91] = 1;
        pixel_data[193][92] = 1;
        pixel_data[193][93] = 6;
        pixel_data[193][94] = 9;
        pixel_data[193][95] = 11;
        pixel_data[193][96] = 9;
        pixel_data[193][97] = 6;
        pixel_data[193][98] = 1;
        pixel_data[193][99] = 1;
        pixel_data[193][100] = 1;
        pixel_data[193][101] = 1;
        pixel_data[193][102] = 1;
        pixel_data[193][103] = 1;
        pixel_data[193][104] = 1;
        pixel_data[193][105] = 1;
        pixel_data[193][106] = 1;
        pixel_data[193][107] = 1;
        pixel_data[193][108] = 1;
        pixel_data[193][109] = 1;
        pixel_data[193][110] = 1;
        pixel_data[193][111] = 1;
        pixel_data[193][112] = 1;
        pixel_data[193][113] = 1;
        pixel_data[193][114] = 1;
        pixel_data[193][115] = 1;
        pixel_data[193][116] = 1;
        pixel_data[193][117] = 1;
        pixel_data[193][118] = 1;
        pixel_data[193][119] = 1;
        pixel_data[193][120] = 1;
        pixel_data[193][121] = 1;
        pixel_data[193][122] = 1;
        pixel_data[193][123] = 1;
        pixel_data[193][124] = 1;
        pixel_data[193][125] = 1;
        pixel_data[193][126] = 1;
        pixel_data[193][127] = 1;
        pixel_data[193][128] = 1;
        pixel_data[193][129] = 1;
        pixel_data[193][130] = 1;
        pixel_data[193][131] = 1;
        pixel_data[193][132] = 1;
        pixel_data[193][133] = 1;
        pixel_data[193][134] = 4;
        pixel_data[193][135] = 4;
        pixel_data[193][136] = 1;
        pixel_data[193][137] = 1;
        pixel_data[193][138] = 1;
        pixel_data[193][139] = 1;
        pixel_data[193][140] = 1;
        pixel_data[193][141] = 1;
        pixel_data[193][142] = 1;
        pixel_data[193][143] = 1;
        pixel_data[193][144] = 1;
        pixel_data[193][145] = 1;
        pixel_data[193][146] = 1;
        pixel_data[193][147] = 1;
        pixel_data[193][148] = 1;
        pixel_data[193][149] = 1;
        pixel_data[193][150] = 1;
        pixel_data[193][151] = 1;
        pixel_data[193][152] = 1;
        pixel_data[193][153] = 1;
        pixel_data[193][154] = 1;
        pixel_data[193][155] = 1;
        pixel_data[193][156] = 1;
        pixel_data[193][157] = 1;
        pixel_data[193][158] = 1;
        pixel_data[193][159] = 1;
        pixel_data[193][160] = 1;
        pixel_data[193][161] = 1;
        pixel_data[193][162] = 1;
        pixel_data[193][163] = 1;
        pixel_data[193][164] = 1;
        pixel_data[193][165] = 1;
        pixel_data[193][166] = 1;
        pixel_data[193][167] = 1;
        pixel_data[193][168] = 1;
        pixel_data[193][169] = 1;
        pixel_data[193][170] = 1;
        pixel_data[193][171] = 1;
        pixel_data[193][172] = 1;
        pixel_data[193][173] = 1;
        pixel_data[193][174] = 1;
        pixel_data[193][175] = 1;
        pixel_data[193][176] = 1;
        pixel_data[193][177] = 1;
        pixel_data[193][178] = 1;
        pixel_data[193][179] = 1;
        pixel_data[193][180] = 1;
        pixel_data[193][181] = 5;
        pixel_data[193][182] = 7;
        pixel_data[193][183] = 9;
        pixel_data[193][184] = 11;
        pixel_data[193][185] = 11;
        pixel_data[193][186] = 0;
        pixel_data[193][187] = 0;
        pixel_data[193][188] = 0;
        pixel_data[193][189] = 0;
        pixel_data[193][190] = 0;
        pixel_data[193][191] = 0;
        pixel_data[193][192] = 0;
        pixel_data[193][193] = 0;
        pixel_data[193][194] = 0;
        pixel_data[193][195] = 0;
        pixel_data[193][196] = 0;
        pixel_data[193][197] = 0;
        pixel_data[193][198] = 0;
        pixel_data[193][199] = 0; // y=193
        pixel_data[194][0] = 0;
        pixel_data[194][1] = 0;
        pixel_data[194][2] = 0;
        pixel_data[194][3] = 0;
        pixel_data[194][4] = 0;
        pixel_data[194][5] = 0;
        pixel_data[194][6] = 0;
        pixel_data[194][7] = 0;
        pixel_data[194][8] = 11;
        pixel_data[194][9] = 11;
        pixel_data[194][10] = 9;
        pixel_data[194][11] = 6;
        pixel_data[194][12] = 1;
        pixel_data[194][13] = 1;
        pixel_data[194][14] = 1;
        pixel_data[194][15] = 1;
        pixel_data[194][16] = 1;
        pixel_data[194][17] = 1;
        pixel_data[194][18] = 4;
        pixel_data[194][19] = 4;
        pixel_data[194][20] = 2;
        pixel_data[194][21] = 1;
        pixel_data[194][22] = 1;
        pixel_data[194][23] = 1;
        pixel_data[194][24] = 1;
        pixel_data[194][25] = 1;
        pixel_data[194][26] = 1;
        pixel_data[194][27] = 1;
        pixel_data[194][28] = 1;
        pixel_data[194][29] = 1;
        pixel_data[194][30] = 1;
        pixel_data[194][31] = 1;
        pixel_data[194][32] = 1;
        pixel_data[194][33] = 1;
        pixel_data[194][34] = 1;
        pixel_data[194][35] = 2;
        pixel_data[194][36] = 4;
        pixel_data[194][37] = 4;
        pixel_data[194][38] = 1;
        pixel_data[194][39] = 1;
        pixel_data[194][40] = 1;
        pixel_data[194][41] = 6;
        pixel_data[194][42] = 8;
        pixel_data[194][43] = 11;
        pixel_data[194][44] = 11;
        pixel_data[194][45] = 0;
        pixel_data[194][46] = 11;
        pixel_data[194][47] = 11;
        pixel_data[194][48] = 8;
        pixel_data[194][49] = 5;
        pixel_data[194][50] = 1;
        pixel_data[194][51] = 1;
        pixel_data[194][52] = 1;
        pixel_data[194][53] = 1;
        pixel_data[194][54] = 1;
        pixel_data[194][55] = 1;
        pixel_data[194][56] = 1;
        pixel_data[194][57] = 1;
        pixel_data[194][58] = 1;
        pixel_data[194][59] = 1;
        pixel_data[194][60] = 1;
        pixel_data[194][61] = 1;
        pixel_data[194][62] = 1;
        pixel_data[194][63] = 1;
        pixel_data[194][64] = 1;
        pixel_data[194][65] = 1;
        pixel_data[194][66] = 1;
        pixel_data[194][67] = 1;
        pixel_data[194][68] = 1;
        pixel_data[194][69] = 1;
        pixel_data[194][70] = 1;
        pixel_data[194][71] = 1;
        pixel_data[194][72] = 1;
        pixel_data[194][73] = 1;
        pixel_data[194][74] = 1;
        pixel_data[194][75] = 1;
        pixel_data[194][76] = 1;
        pixel_data[194][77] = 1;
        pixel_data[194][78] = 1;
        pixel_data[194][79] = 1;
        pixel_data[194][80] = 1;
        pixel_data[194][81] = 1;
        pixel_data[194][82] = 1;
        pixel_data[194][83] = 1;
        pixel_data[194][84] = 1;
        pixel_data[194][85] = 1;
        pixel_data[194][86] = 1;
        pixel_data[194][87] = 1;
        pixel_data[194][88] = 1;
        pixel_data[194][89] = 1;
        pixel_data[194][90] = 1;
        pixel_data[194][91] = 1;
        pixel_data[194][92] = 6;
        pixel_data[194][93] = 9;
        pixel_data[194][94] = 11;
        pixel_data[194][95] = 11;
        pixel_data[194][96] = 11;
        pixel_data[194][97] = 9;
        pixel_data[194][98] = 7;
        pixel_data[194][99] = 1;
        pixel_data[194][100] = 1;
        pixel_data[194][101] = 1;
        pixel_data[194][102] = 1;
        pixel_data[194][103] = 1;
        pixel_data[194][104] = 1;
        pixel_data[194][105] = 1;
        pixel_data[194][106] = 1;
        pixel_data[194][107] = 1;
        pixel_data[194][108] = 1;
        pixel_data[194][109] = 1;
        pixel_data[194][110] = 1;
        pixel_data[194][111] = 1;
        pixel_data[194][112] = 1;
        pixel_data[194][113] = 1;
        pixel_data[194][114] = 1;
        pixel_data[194][115] = 1;
        pixel_data[194][116] = 1;
        pixel_data[194][117] = 1;
        pixel_data[194][118] = 1;
        pixel_data[194][119] = 1;
        pixel_data[194][120] = 1;
        pixel_data[194][121] = 1;
        pixel_data[194][122] = 1;
        pixel_data[194][123] = 1;
        pixel_data[194][124] = 1;
        pixel_data[194][125] = 1;
        pixel_data[194][126] = 1;
        pixel_data[194][127] = 1;
        pixel_data[194][128] = 1;
        pixel_data[194][129] = 1;
        pixel_data[194][130] = 1;
        pixel_data[194][131] = 1;
        pixel_data[194][132] = 6;
        pixel_data[194][133] = 8;
        pixel_data[194][134] = 11;
        pixel_data[194][135] = 11;
        pixel_data[194][136] = 9;
        pixel_data[194][137] = 7;
        pixel_data[194][138] = 2;
        pixel_data[194][139] = 1;
        pixel_data[194][140] = 1;
        pixel_data[194][141] = 1;
        pixel_data[194][142] = 1;
        pixel_data[194][143] = 1;
        pixel_data[194][144] = 1;
        pixel_data[194][145] = 1;
        pixel_data[194][146] = 1;
        pixel_data[194][147] = 1;
        pixel_data[194][148] = 1;
        pixel_data[194][149] = 1;
        pixel_data[194][150] = 1;
        pixel_data[194][151] = 1;
        pixel_data[194][152] = 1;
        pixel_data[194][153] = 1;
        pixel_data[194][154] = 1;
        pixel_data[194][155] = 1;
        pixel_data[194][156] = 1;
        pixel_data[194][157] = 1;
        pixel_data[194][158] = 1;
        pixel_data[194][159] = 1;
        pixel_data[194][160] = 1;
        pixel_data[194][161] = 1;
        pixel_data[194][162] = 1;
        pixel_data[194][163] = 1;
        pixel_data[194][164] = 1;
        pixel_data[194][165] = 1;
        pixel_data[194][166] = 1;
        pixel_data[194][167] = 1;
        pixel_data[194][168] = 1;
        pixel_data[194][169] = 1;
        pixel_data[194][170] = 1;
        pixel_data[194][171] = 1;
        pixel_data[194][172] = 1;
        pixel_data[194][173] = 1;
        pixel_data[194][174] = 1;
        pixel_data[194][175] = 1;
        pixel_data[194][176] = 1;
        pixel_data[194][177] = 1;
        pixel_data[194][178] = 4;
        pixel_data[194][179] = 6;
        pixel_data[194][180] = 8;
        pixel_data[194][181] = 9;
        pixel_data[194][182] = 11;
        pixel_data[194][183] = 11;
        pixel_data[194][184] = 0;
        pixel_data[194][185] = 0;
        pixel_data[194][186] = 0;
        pixel_data[194][187] = 0;
        pixel_data[194][188] = 0;
        pixel_data[194][189] = 0;
        pixel_data[194][190] = 0;
        pixel_data[194][191] = 0;
        pixel_data[194][192] = 0;
        pixel_data[194][193] = 0;
        pixel_data[194][194] = 0;
        pixel_data[194][195] = 0;
        pixel_data[194][196] = 0;
        pixel_data[194][197] = 0;
        pixel_data[194][198] = 0;
        pixel_data[194][199] = 0; // y=194
        pixel_data[195][0] = 0;
        pixel_data[195][1] = 0;
        pixel_data[195][2] = 0;
        pixel_data[195][3] = 0;
        pixel_data[195][4] = 0;
        pixel_data[195][5] = 0;
        pixel_data[195][6] = 0;
        pixel_data[195][7] = 0;
        pixel_data[195][8] = 0;
        pixel_data[195][9] = 11;
        pixel_data[195][10] = 11;
        pixel_data[195][11] = 9;
        pixel_data[195][12] = 8;
        pixel_data[195][13] = 5;
        pixel_data[195][14] = 1;
        pixel_data[195][15] = 1;
        pixel_data[195][16] = 1;
        pixel_data[195][17] = 1;
        pixel_data[195][18] = 1;
        pixel_data[195][19] = 4;
        pixel_data[195][20] = 4;
        pixel_data[195][21] = 2;
        pixel_data[195][22] = 1;
        pixel_data[195][23] = 1;
        pixel_data[195][24] = 1;
        pixel_data[195][25] = 1;
        pixel_data[195][26] = 1;
        pixel_data[195][27] = 1;
        pixel_data[195][28] = 1;
        pixel_data[195][29] = 1;
        pixel_data[195][30] = 1;
        pixel_data[195][31] = 1;
        pixel_data[195][32] = 1;
        pixel_data[195][33] = 1;
        pixel_data[195][34] = 2;
        pixel_data[195][35] = 4;
        pixel_data[195][36] = 4;
        pixel_data[195][37] = 1;
        pixel_data[195][38] = 1;
        pixel_data[195][39] = 2;
        pixel_data[195][40] = 7;
        pixel_data[195][41] = 9;
        pixel_data[195][42] = 11;
        pixel_data[195][43] = 11;
        pixel_data[195][44] = 0;
        pixel_data[195][45] = 0;
        pixel_data[195][46] = 0;
        pixel_data[195][47] = 10;
        pixel_data[195][48] = 11;
        pixel_data[195][49] = 9;
        pixel_data[195][50] = 8;
        pixel_data[195][51] = 4;
        pixel_data[195][52] = 1;
        pixel_data[195][53] = 1;
        pixel_data[195][54] = 1;
        pixel_data[195][55] = 1;
        pixel_data[195][56] = 1;
        pixel_data[195][57] = 1;
        pixel_data[195][58] = 1;
        pixel_data[195][59] = 1;
        pixel_data[195][60] = 1;
        pixel_data[195][61] = 1;
        pixel_data[195][62] = 1;
        pixel_data[195][63] = 1;
        pixel_data[195][64] = 1;
        pixel_data[195][65] = 1;
        pixel_data[195][66] = 1;
        pixel_data[195][67] = 1;
        pixel_data[195][68] = 1;
        pixel_data[195][69] = 1;
        pixel_data[195][70] = 1;
        pixel_data[195][71] = 1;
        pixel_data[195][72] = 1;
        pixel_data[195][73] = 1;
        pixel_data[195][74] = 1;
        pixel_data[195][75] = 1;
        pixel_data[195][76] = 1;
        pixel_data[195][77] = 1;
        pixel_data[195][78] = 1;
        pixel_data[195][79] = 1;
        pixel_data[195][80] = 1;
        pixel_data[195][81] = 1;
        pixel_data[195][82] = 1;
        pixel_data[195][83] = 1;
        pixel_data[195][84] = 1;
        pixel_data[195][85] = 1;
        pixel_data[195][86] = 1;
        pixel_data[195][87] = 1;
        pixel_data[195][88] = 1;
        pixel_data[195][89] = 2;
        pixel_data[195][90] = 6;
        pixel_data[195][91] = 9;
        pixel_data[195][92] = 11;
        pixel_data[195][93] = 11;
        pixel_data[195][94] = 0;
        pixel_data[195][95] = 0;
        pixel_data[195][96] = 0;
        pixel_data[195][97] = 11;
        pixel_data[195][98] = 11;
        pixel_data[195][99] = 9;
        pixel_data[195][100] = 7;
        pixel_data[195][101] = 2;
        pixel_data[195][102] = 1;
        pixel_data[195][103] = 1;
        pixel_data[195][104] = 1;
        pixel_data[195][105] = 1;
        pixel_data[195][106] = 1;
        pixel_data[195][107] = 1;
        pixel_data[195][108] = 1;
        pixel_data[195][109] = 1;
        pixel_data[195][110] = 1;
        pixel_data[195][111] = 1;
        pixel_data[195][112] = 1;
        pixel_data[195][113] = 1;
        pixel_data[195][114] = 1;
        pixel_data[195][115] = 1;
        pixel_data[195][116] = 1;
        pixel_data[195][117] = 1;
        pixel_data[195][118] = 1;
        pixel_data[195][119] = 1;
        pixel_data[195][120] = 1;
        pixel_data[195][121] = 1;
        pixel_data[195][122] = 1;
        pixel_data[195][123] = 1;
        pixel_data[195][124] = 1;
        pixel_data[195][125] = 1;
        pixel_data[195][126] = 1;
        pixel_data[195][127] = 1;
        pixel_data[195][128] = 1;
        pixel_data[195][129] = 1;
        pixel_data[195][130] = 5;
        pixel_data[195][131] = 8;
        pixel_data[195][132] = 11;
        pixel_data[195][133] = 11;
        pixel_data[195][134] = 0;
        pixel_data[195][135] = 0;
        pixel_data[195][136] = 11;
        pixel_data[195][137] = 11;
        pixel_data[195][138] = 9;
        pixel_data[195][139] = 7;
        pixel_data[195][140] = 2;
        pixel_data[195][141] = 1;
        pixel_data[195][142] = 1;
        pixel_data[195][143] = 1;
        pixel_data[195][144] = 1;
        pixel_data[195][145] = 1;
        pixel_data[195][146] = 1;
        pixel_data[195][147] = 1;
        pixel_data[195][148] = 1;
        pixel_data[195][149] = 1;
        pixel_data[195][150] = 1;
        pixel_data[195][151] = 1;
        pixel_data[195][152] = 1;
        pixel_data[195][153] = 1;
        pixel_data[195][154] = 1;
        pixel_data[195][155] = 1;
        pixel_data[195][156] = 1;
        pixel_data[195][157] = 1;
        pixel_data[195][158] = 1;
        pixel_data[195][159] = 1;
        pixel_data[195][160] = 1;
        pixel_data[195][161] = 1;
        pixel_data[195][162] = 1;
        pixel_data[195][163] = 1;
        pixel_data[195][164] = 1;
        pixel_data[195][165] = 1;
        pixel_data[195][166] = 1;
        pixel_data[195][167] = 1;
        pixel_data[195][168] = 1;
        pixel_data[195][169] = 1;
        pixel_data[195][170] = 1;
        pixel_data[195][171] = 1;
        pixel_data[195][172] = 1;
        pixel_data[195][173] = 4;
        pixel_data[195][174] = 6;
        pixel_data[195][175] = 8;
        pixel_data[195][176] = 9;
        pixel_data[195][177] = 11;
        pixel_data[195][178] = 11;
        pixel_data[195][179] = 10;
        pixel_data[195][180] = 0;
        pixel_data[195][181] = 0;
        pixel_data[195][182] = 0;
        pixel_data[195][183] = 0;
        pixel_data[195][184] = 0;
        pixel_data[195][185] = 0;
        pixel_data[195][186] = 0;
        pixel_data[195][187] = 0;
        pixel_data[195][188] = 0;
        pixel_data[195][189] = 0;
        pixel_data[195][190] = 0;
        pixel_data[195][191] = 0;
        pixel_data[195][192] = 0;
        pixel_data[195][193] = 0;
        pixel_data[195][194] = 0;
        pixel_data[195][195] = 0;
        pixel_data[195][196] = 0;
        pixel_data[195][197] = 0;
        pixel_data[195][198] = 0;
        pixel_data[195][199] = 0; // y=195
        pixel_data[196][0] = 0;
        pixel_data[196][1] = 0;
        pixel_data[196][2] = 0;
        pixel_data[196][3] = 0;
        pixel_data[196][4] = 0;
        pixel_data[196][5] = 0;
        pixel_data[196][6] = 0;
        pixel_data[196][7] = 0;
        pixel_data[196][8] = 0;
        pixel_data[196][9] = 0;
        pixel_data[196][10] = 0;
        pixel_data[196][11] = 11;
        pixel_data[196][12] = 11;
        pixel_data[196][13] = 9;
        pixel_data[196][14] = 6;
        pixel_data[196][15] = 1;
        pixel_data[196][16] = 1;
        pixel_data[196][17] = 1;
        pixel_data[196][18] = 1;
        pixel_data[196][19] = 2;
        pixel_data[196][20] = 4;
        pixel_data[196][21] = 4;
        pixel_data[196][22] = 1;
        pixel_data[196][23] = 1;
        pixel_data[196][24] = 1;
        pixel_data[196][25] = 1;
        pixel_data[196][26] = 1;
        pixel_data[196][27] = 1;
        pixel_data[196][28] = 1;
        pixel_data[196][29] = 1;
        pixel_data[196][30] = 1;
        pixel_data[196][31] = 1;
        pixel_data[196][32] = 1;
        pixel_data[196][33] = 2;
        pixel_data[196][34] = 4;
        pixel_data[196][35] = 4;
        pixel_data[196][36] = 1;
        pixel_data[196][37] = 1;
        pixel_data[196][38] = 5;
        pixel_data[196][39] = 8;
        pixel_data[196][40] = 9;
        pixel_data[196][41] = 11;
        pixel_data[196][42] = 11;
        pixel_data[196][43] = 0;
        pixel_data[196][44] = 0;
        pixel_data[196][45] = 0;
        pixel_data[196][46] = 0;
        pixel_data[196][47] = 0;
        pixel_data[196][48] = 0;
        pixel_data[196][49] = 11;
        pixel_data[196][50] = 11;
        pixel_data[196][51] = 9;
        pixel_data[196][52] = 7;
        pixel_data[196][53] = 4;
        pixel_data[196][54] = 1;
        pixel_data[196][55] = 1;
        pixel_data[196][56] = 1;
        pixel_data[196][57] = 1;
        pixel_data[196][58] = 1;
        pixel_data[196][59] = 1;
        pixel_data[196][60] = 1;
        pixel_data[196][61] = 1;
        pixel_data[196][62] = 1;
        pixel_data[196][63] = 1;
        pixel_data[196][64] = 1;
        pixel_data[196][65] = 1;
        pixel_data[196][66] = 1;
        pixel_data[196][67] = 1;
        pixel_data[196][68] = 1;
        pixel_data[196][69] = 1;
        pixel_data[196][70] = 1;
        pixel_data[196][71] = 1;
        pixel_data[196][72] = 1;
        pixel_data[196][73] = 1;
        pixel_data[196][74] = 1;
        pixel_data[196][75] = 1;
        pixel_data[196][76] = 1;
        pixel_data[196][77] = 1;
        pixel_data[196][78] = 1;
        pixel_data[196][79] = 1;
        pixel_data[196][80] = 1;
        pixel_data[196][81] = 1;
        pixel_data[196][82] = 1;
        pixel_data[196][83] = 1;
        pixel_data[196][84] = 1;
        pixel_data[196][85] = 1;
        pixel_data[196][86] = 1;
        pixel_data[196][87] = 1;
        pixel_data[196][88] = 6;
        pixel_data[196][89] = 8;
        pixel_data[196][90] = 11;
        pixel_data[196][91] = 11;
        pixel_data[196][92] = 13;
        pixel_data[196][93] = 0;
        pixel_data[196][94] = 0;
        pixel_data[196][95] = 0;
        pixel_data[196][96] = 0;
        pixel_data[196][97] = 0;
        pixel_data[196][98] = 0;
        pixel_data[196][99] = 11;
        pixel_data[196][100] = 11;
        pixel_data[196][101] = 9;
        pixel_data[196][102] = 7;
        pixel_data[196][103] = 5;
        pixel_data[196][104] = 1;
        pixel_data[196][105] = 1;
        pixel_data[196][106] = 1;
        pixel_data[196][107] = 1;
        pixel_data[196][108] = 1;
        pixel_data[196][109] = 1;
        pixel_data[196][110] = 1;
        pixel_data[196][111] = 1;
        pixel_data[196][112] = 1;
        pixel_data[196][113] = 1;
        pixel_data[196][114] = 1;
        pixel_data[196][115] = 1;
        pixel_data[196][116] = 1;
        pixel_data[196][117] = 1;
        pixel_data[196][118] = 1;
        pixel_data[196][119] = 1;
        pixel_data[196][120] = 1;
        pixel_data[196][121] = 1;
        pixel_data[196][122] = 1;
        pixel_data[196][123] = 1;
        pixel_data[196][124] = 1;
        pixel_data[196][125] = 1;
        pixel_data[196][126] = 1;
        pixel_data[196][127] = 1;
        pixel_data[196][128] = 1;
        pixel_data[196][129] = 6;
        pixel_data[196][130] = 8;
        pixel_data[196][131] = 11;
        pixel_data[196][132] = 11;
        pixel_data[196][133] = 0;
        pixel_data[196][134] = 0;
        pixel_data[196][135] = 0;
        pixel_data[196][136] = 0;
        pixel_data[196][137] = 13;
        pixel_data[196][138] = 11;
        pixel_data[196][139] = 11;
        pixel_data[196][140] = 8;
        pixel_data[196][141] = 5;
        pixel_data[196][142] = 1;
        pixel_data[196][143] = 1;
        pixel_data[196][144] = 1;
        pixel_data[196][145] = 1;
        pixel_data[196][146] = 1;
        pixel_data[196][147] = 1;
        pixel_data[196][148] = 1;
        pixel_data[196][149] = 1;
        pixel_data[196][150] = 1;
        pixel_data[196][151] = 1;
        pixel_data[196][152] = 1;
        pixel_data[196][153] = 1;
        pixel_data[196][154] = 1;
        pixel_data[196][155] = 1;
        pixel_data[196][156] = 1;
        pixel_data[196][157] = 1;
        pixel_data[196][158] = 1;
        pixel_data[196][159] = 1;
        pixel_data[196][160] = 1;
        pixel_data[196][161] = 1;
        pixel_data[196][162] = 1;
        pixel_data[196][163] = 1;
        pixel_data[196][164] = 1;
        pixel_data[196][165] = 1;
        pixel_data[196][166] = 1;
        pixel_data[196][167] = 1;
        pixel_data[196][168] = 1;
        pixel_data[196][169] = 1;
        pixel_data[196][170] = 5;
        pixel_data[196][171] = 7;
        pixel_data[196][172] = 9;
        pixel_data[196][173] = 11;
        pixel_data[196][174] = 11;
        pixel_data[196][175] = 11;
        pixel_data[196][176] = 0;
        pixel_data[196][177] = 0;
        pixel_data[196][178] = 0;
        pixel_data[196][179] = 0;
        pixel_data[196][180] = 0;
        pixel_data[196][181] = 0;
        pixel_data[196][182] = 0;
        pixel_data[196][183] = 0;
        pixel_data[196][184] = 0;
        pixel_data[196][185] = 0;
        pixel_data[196][186] = 0;
        pixel_data[196][187] = 0;
        pixel_data[196][188] = 0;
        pixel_data[196][189] = 0;
        pixel_data[196][190] = 0;
        pixel_data[196][191] = 0;
        pixel_data[196][192] = 0;
        pixel_data[196][193] = 0;
        pixel_data[196][194] = 0;
        pixel_data[196][195] = 0;
        pixel_data[196][196] = 0;
        pixel_data[196][197] = 0;
        pixel_data[196][198] = 0;
        pixel_data[196][199] = 0; // y=196
        pixel_data[197][0] = 0;
        pixel_data[197][1] = 0;
        pixel_data[197][2] = 0;
        pixel_data[197][3] = 0;
        pixel_data[197][4] = 0;
        pixel_data[197][5] = 0;
        pixel_data[197][6] = 0;
        pixel_data[197][7] = 0;
        pixel_data[197][8] = 0;
        pixel_data[197][9] = 0;
        pixel_data[197][10] = 0;
        pixel_data[197][11] = 0;
        pixel_data[197][12] = 0;
        pixel_data[197][13] = 11;
        pixel_data[197][14] = 11;
        pixel_data[197][15] = 9;
        pixel_data[197][16] = 8;
        pixel_data[197][17] = 6;
        pixel_data[197][18] = 2;
        pixel_data[197][19] = 1;
        pixel_data[197][20] = 1;
        pixel_data[197][21] = 4;
        pixel_data[197][22] = 4;
        pixel_data[197][23] = 4;
        pixel_data[197][24] = 2;
        pixel_data[197][25] = 2;
        pixel_data[197][26] = 2;
        pixel_data[197][27] = 2;
        pixel_data[197][28] = 2;
        pixel_data[197][29] = 2;
        pixel_data[197][30] = 4;
        pixel_data[197][31] = 4;
        pixel_data[197][32] = 4;
        pixel_data[197][33] = 4;
        pixel_data[197][34] = 1;
        pixel_data[197][35] = 5;
        pixel_data[197][36] = 7;
        pixel_data[197][37] = 9;
        pixel_data[197][38] = 11;
        pixel_data[197][39] = 11;
        pixel_data[197][40] = 11;
        pixel_data[197][41] = 0;
        pixel_data[197][42] = 0;
        pixel_data[197][43] = 0;
        pixel_data[197][44] = 0;
        pixel_data[197][45] = 0;
        pixel_data[197][46] = 0;
        pixel_data[197][47] = 0;
        pixel_data[197][48] = 0;
        pixel_data[197][49] = 0;
        pixel_data[197][50] = 0;
        pixel_data[197][51] = 11;
        pixel_data[197][52] = 11;
        pixel_data[197][53] = 9;
        pixel_data[197][54] = 8;
        pixel_data[197][55] = 5;
        pixel_data[197][56] = 1;
        pixel_data[197][57] = 1;
        pixel_data[197][58] = 1;
        pixel_data[197][59] = 1;
        pixel_data[197][60] = 1;
        pixel_data[197][61] = 1;
        pixel_data[197][62] = 1;
        pixel_data[197][63] = 1;
        pixel_data[197][64] = 1;
        pixel_data[197][65] = 1;
        pixel_data[197][66] = 1;
        pixel_data[197][67] = 1;
        pixel_data[197][68] = 1;
        pixel_data[197][69] = 1;
        pixel_data[197][70] = 1;
        pixel_data[197][71] = 1;
        pixel_data[197][72] = 1;
        pixel_data[197][73] = 1;
        pixel_data[197][74] = 1;
        pixel_data[197][75] = 1;
        pixel_data[197][76] = 1;
        pixel_data[197][77] = 1;
        pixel_data[197][78] = 1;
        pixel_data[197][79] = 1;
        pixel_data[197][80] = 1;
        pixel_data[197][81] = 1;
        pixel_data[197][82] = 1;
        pixel_data[197][83] = 1;
        pixel_data[197][84] = 1;
        pixel_data[197][85] = 1;
        pixel_data[197][86] = 6;
        pixel_data[197][87] = 8;
        pixel_data[197][88] = 11;
        pixel_data[197][89] = 11;
        pixel_data[197][90] = 11;
        pixel_data[197][91] = 0;
        pixel_data[197][92] = 0;
        pixel_data[197][93] = 0;
        pixel_data[197][94] = 0;
        pixel_data[197][95] = 0;
        pixel_data[197][96] = 0;
        pixel_data[197][97] = 0;
        pixel_data[197][98] = 0;
        pixel_data[197][99] = 0;
        pixel_data[197][100] = 0;
        pixel_data[197][101] = 10;
        pixel_data[197][102] = 11;
        pixel_data[197][103] = 11;
        pixel_data[197][104] = 9;
        pixel_data[197][105] = 8;
        pixel_data[197][106] = 7;
        pixel_data[197][107] = 5;
        pixel_data[197][108] = 1;
        pixel_data[197][109] = 1;
        pixel_data[197][110] = 1;
        pixel_data[197][111] = 1;
        pixel_data[197][112] = 1;
        pixel_data[197][113] = 1;
        pixel_data[197][114] = 1;
        pixel_data[197][115] = 1;
        pixel_data[197][116] = 1;
        pixel_data[197][117] = 1;
        pixel_data[197][118] = 1;
        pixel_data[197][119] = 1;
        pixel_data[197][120] = 1;
        pixel_data[197][121] = 1;
        pixel_data[197][122] = 1;
        pixel_data[197][123] = 1;
        pixel_data[197][124] = 1;
        pixel_data[197][125] = 4;
        pixel_data[197][126] = 6;
        pixel_data[197][127] = 8;
        pixel_data[197][128] = 9;
        pixel_data[197][129] = 11;
        pixel_data[197][130] = 11;
        pixel_data[197][131] = 13;
        pixel_data[197][132] = 0;
        pixel_data[197][133] = 0;
        pixel_data[197][134] = 0;
        pixel_data[197][135] = 0;
        pixel_data[197][136] = 0;
        pixel_data[197][137] = 0;
        pixel_data[197][138] = 0;
        pixel_data[197][139] = 9;
        pixel_data[197][140] = 11;
        pixel_data[197][141] = 9;
        pixel_data[197][142] = 8;
        pixel_data[197][143] = 7;
        pixel_data[197][144] = 5;
        pixel_data[197][145] = 1;
        pixel_data[197][146] = 1;
        pixel_data[197][147] = 1;
        pixel_data[197][148] = 1;
        pixel_data[197][149] = 1;
        pixel_data[197][150] = 1;
        pixel_data[197][151] = 1;
        pixel_data[197][152] = 1;
        pixel_data[197][153] = 1;
        pixel_data[197][154] = 1;
        pixel_data[197][155] = 1;
        pixel_data[197][156] = 1;
        pixel_data[197][157] = 1;
        pixel_data[197][158] = 1;
        pixel_data[197][159] = 1;
        pixel_data[197][160] = 1;
        pixel_data[197][161] = 1;
        pixel_data[197][162] = 1;
        pixel_data[197][163] = 1;
        pixel_data[197][164] = 1;
        pixel_data[197][165] = 4;
        pixel_data[197][166] = 6;
        pixel_data[197][167] = 7;
        pixel_data[197][168] = 8;
        pixel_data[197][169] = 9;
        pixel_data[197][170] = 11;
        pixel_data[197][171] = 11;
        pixel_data[197][172] = 11;
        pixel_data[197][173] = 0;
        pixel_data[197][174] = 0;
        pixel_data[197][175] = 0;
        pixel_data[197][176] = 0;
        pixel_data[197][177] = 0;
        pixel_data[197][178] = 0;
        pixel_data[197][179] = 0;
        pixel_data[197][180] = 0;
        pixel_data[197][181] = 0;
        pixel_data[197][182] = 0;
        pixel_data[197][183] = 0;
        pixel_data[197][184] = 0;
        pixel_data[197][185] = 0;
        pixel_data[197][186] = 0;
        pixel_data[197][187] = 0;
        pixel_data[197][188] = 0;
        pixel_data[197][189] = 0;
        pixel_data[197][190] = 0;
        pixel_data[197][191] = 0;
        pixel_data[197][192] = 0;
        pixel_data[197][193] = 0;
        pixel_data[197][194] = 0;
        pixel_data[197][195] = 0;
        pixel_data[197][196] = 0;
        pixel_data[197][197] = 0;
        pixel_data[197][198] = 0;
        pixel_data[197][199] = 0; // y=197
        pixel_data[198][0] = 0;
        pixel_data[198][1] = 0;
        pixel_data[198][2] = 0;
        pixel_data[198][3] = 0;
        pixel_data[198][4] = 0;
        pixel_data[198][5] = 0;
        pixel_data[198][6] = 0;
        pixel_data[198][7] = 0;
        pixel_data[198][8] = 0;
        pixel_data[198][9] = 0;
        pixel_data[198][10] = 0;
        pixel_data[198][11] = 0;
        pixel_data[198][12] = 0;
        pixel_data[198][13] = 0;
        pixel_data[198][14] = 0;
        pixel_data[198][15] = 0;
        pixel_data[198][16] = 0;
        pixel_data[198][17] = 11;
        pixel_data[198][18] = 11;
        pixel_data[198][19] = 11;
        pixel_data[198][20] = 11;
        pixel_data[198][21] = 9;
        pixel_data[198][22] = 9;
        pixel_data[198][23] = 9;
        pixel_data[198][24] = 8;
        pixel_data[198][25] = 8;
        pixel_data[198][26] = 8;
        pixel_data[198][27] = 8;
        pixel_data[198][28] = 8;
        pixel_data[198][29] = 8;
        pixel_data[198][30] = 8;
        pixel_data[198][31] = 8;
        pixel_data[198][32] = 9;
        pixel_data[198][33] = 11;
        pixel_data[198][34] = 11;
        pixel_data[198][35] = 11;
        pixel_data[198][36] = 13;
        pixel_data[198][37] = 0;
        pixel_data[198][38] = 0;
        pixel_data[198][39] = 0;
        pixel_data[198][40] = 0;
        pixel_data[198][41] = 0;
        pixel_data[198][42] = 0;
        pixel_data[198][43] = 0;
        pixel_data[198][44] = 0;
        pixel_data[198][45] = 0;
        pixel_data[198][46] = 0;
        pixel_data[198][47] = 0;
        pixel_data[198][48] = 0;
        pixel_data[198][49] = 0;
        pixel_data[198][50] = 0;
        pixel_data[198][51] = 0;
        pixel_data[198][52] = 0;
        pixel_data[198][53] = 0;
        pixel_data[198][54] = 0;
        pixel_data[198][55] = 11;
        pixel_data[198][56] = 11;
        pixel_data[198][57] = 11;
        pixel_data[198][58] = 9;
        pixel_data[198][59] = 8;
        pixel_data[198][60] = 7;
        pixel_data[198][61] = 6;
        pixel_data[198][62] = 5;
        pixel_data[198][63] = 2;
        pixel_data[198][64] = 1;
        pixel_data[198][65] = 1;
        pixel_data[198][66] = 1;
        pixel_data[198][67] = 1;
        pixel_data[198][68] = 1;
        pixel_data[198][69] = 1;
        pixel_data[198][70] = 1;
        pixel_data[198][71] = 1;
        pixel_data[198][72] = 1;
        pixel_data[198][73] = 1;
        pixel_data[198][74] = 1;
        pixel_data[198][75] = 1;
        pixel_data[198][76] = 1;
        pixel_data[198][77] = 1;
        pixel_data[198][78] = 1;
        pixel_data[198][79] = 1;
        pixel_data[198][80] = 1;
        pixel_data[198][81] = 4;
        pixel_data[198][82] = 6;
        pixel_data[198][83] = 7;
        pixel_data[198][84] = 9;
        pixel_data[198][85] = 11;
        pixel_data[198][86] = 11;
        pixel_data[198][87] = 11;
        pixel_data[198][88] = 0;
        pixel_data[198][89] = 0;
        pixel_data[198][90] = 0;
        pixel_data[198][91] = 0;
        pixel_data[198][92] = 0;
        pixel_data[198][93] = 0;
        pixel_data[198][94] = 0;
        pixel_data[198][95] = 0;
        pixel_data[198][96] = 0;
        pixel_data[198][97] = 0;
        pixel_data[198][98] = 0;
        pixel_data[198][99] = 0;
        pixel_data[198][100] = 0;
        pixel_data[198][101] = 0;
        pixel_data[198][102] = 0;
        pixel_data[198][103] = 0;
        pixel_data[198][104] = 0;
        pixel_data[198][105] = 0;
        pixel_data[198][106] = 0;
        pixel_data[198][107] = 11;
        pixel_data[198][108] = 11;
        pixel_data[198][109] = 11;
        pixel_data[198][110] = 11;
        pixel_data[198][111] = 11;
        pixel_data[198][112] = 11;
        pixel_data[198][113] = 11;
        pixel_data[198][114] = 11;
        pixel_data[198][115] = 11;
        pixel_data[198][116] = 9;
        pixel_data[198][117] = 9;
        pixel_data[198][118] = 9;
        pixel_data[198][119] = 9;
        pixel_data[198][120] = 9;
        pixel_data[198][121] = 9;
        pixel_data[198][122] = 11;
        pixel_data[198][123] = 11;
        pixel_data[198][124] = 11;
        pixel_data[198][125] = 11;
        pixel_data[198][126] = 0;
        pixel_data[198][127] = 0;
        pixel_data[198][128] = 0;
        pixel_data[198][129] = 0;
        pixel_data[198][130] = 0;
        pixel_data[198][131] = 0;
        pixel_data[198][132] = 0;
        pixel_data[198][133] = 0;
        pixel_data[198][134] = 0;
        pixel_data[198][135] = 0;
        pixel_data[198][136] = 0;
        pixel_data[198][137] = 0;
        pixel_data[198][138] = 0;
        pixel_data[198][139] = 0;
        pixel_data[198][140] = 0;
        pixel_data[198][141] = 0;
        pixel_data[198][142] = 0;
        pixel_data[198][143] = 0;
        pixel_data[198][144] = 0;
        pixel_data[198][145] = 10;
        pixel_data[198][146] = 11;
        pixel_data[198][147] = 11;
        pixel_data[198][148] = 11;
        pixel_data[198][149] = 11;
        pixel_data[198][150] = 11;
        pixel_data[198][151] = 11;
        pixel_data[198][152] = 11;
        pixel_data[198][153] = 11;
        pixel_data[198][154] = 11;
        pixel_data[198][155] = 11;
        pixel_data[198][156] = 11;
        pixel_data[198][157] = 11;
        pixel_data[198][158] = 11;
        pixel_data[198][159] = 11;
        pixel_data[198][160] = 11;
        pixel_data[198][161] = 11;
        pixel_data[198][162] = 11;
        pixel_data[198][163] = 11;
        pixel_data[198][164] = 11;
        pixel_data[198][165] = 0;
        pixel_data[198][166] = 0;
        pixel_data[198][167] = 0;
        pixel_data[198][168] = 0;
        pixel_data[198][169] = 0;
        pixel_data[198][170] = 0;
        pixel_data[198][171] = 0;
        pixel_data[198][172] = 0;
        pixel_data[198][173] = 0;
        pixel_data[198][174] = 0;
        pixel_data[198][175] = 0;
        pixel_data[198][176] = 0;
        pixel_data[198][177] = 0;
        pixel_data[198][178] = 0;
        pixel_data[198][179] = 0;
        pixel_data[198][180] = 0;
        pixel_data[198][181] = 0;
        pixel_data[198][182] = 0;
        pixel_data[198][183] = 0;
        pixel_data[198][184] = 0;
        pixel_data[198][185] = 0;
        pixel_data[198][186] = 0;
        pixel_data[198][187] = 0;
        pixel_data[198][188] = 0;
        pixel_data[198][189] = 0;
        pixel_data[198][190] = 0;
        pixel_data[198][191] = 0;
        pixel_data[198][192] = 0;
        pixel_data[198][193] = 0;
        pixel_data[198][194] = 0;
        pixel_data[198][195] = 0;
        pixel_data[198][196] = 0;
        pixel_data[198][197] = 0;
        pixel_data[198][198] = 0;
        pixel_data[198][199] = 0; // y=198
        pixel_data[199][0] = 0;
        pixel_data[199][1] = 0;
        pixel_data[199][2] = 0;
        pixel_data[199][3] = 0;
        pixel_data[199][4] = 0;
        pixel_data[199][5] = 0;
        pixel_data[199][6] = 0;
        pixel_data[199][7] = 0;
        pixel_data[199][8] = 0;
        pixel_data[199][9] = 0;
        pixel_data[199][10] = 0;
        pixel_data[199][11] = 0;
        pixel_data[199][12] = 0;
        pixel_data[199][13] = 0;
        pixel_data[199][14] = 0;
        pixel_data[199][15] = 0;
        pixel_data[199][16] = 0;
        pixel_data[199][17] = 0;
        pixel_data[199][18] = 0;
        pixel_data[199][19] = 0;
        pixel_data[199][20] = 0;
        pixel_data[199][21] = 0;
        pixel_data[199][22] = 0;
        pixel_data[199][23] = 0;
        pixel_data[199][24] = 0;
        pixel_data[199][25] = 0;
        pixel_data[199][26] = 0;
        pixel_data[199][27] = 0;
        pixel_data[199][28] = 0;
        pixel_data[199][29] = 0;
        pixel_data[199][30] = 0;
        pixel_data[199][31] = 0;
        pixel_data[199][32] = 0;
        pixel_data[199][33] = 0;
        pixel_data[199][34] = 0;
        pixel_data[199][35] = 0;
        pixel_data[199][36] = 0;
        pixel_data[199][37] = 0;
        pixel_data[199][38] = 0;
        pixel_data[199][39] = 0;
        pixel_data[199][40] = 0;
        pixel_data[199][41] = 0;
        pixel_data[199][42] = 0;
        pixel_data[199][43] = 0;
        pixel_data[199][44] = 0;
        pixel_data[199][45] = 0;
        pixel_data[199][46] = 0;
        pixel_data[199][47] = 0;
        pixel_data[199][48] = 0;
        pixel_data[199][49] = 0;
        pixel_data[199][50] = 0;
        pixel_data[199][51] = 0;
        pixel_data[199][52] = 0;
        pixel_data[199][53] = 0;
        pixel_data[199][54] = 0;
        pixel_data[199][55] = 0;
        pixel_data[199][56] = 0;
        pixel_data[199][57] = 0;
        pixel_data[199][58] = 0;
        pixel_data[199][59] = 0;
        pixel_data[199][60] = 11;
        pixel_data[199][61] = 11;
        pixel_data[199][62] = 11;
        pixel_data[199][63] = 11;
        pixel_data[199][64] = 11;
        pixel_data[199][65] = 11;
        pixel_data[199][66] = 11;
        pixel_data[199][67] = 11;
        pixel_data[199][68] = 9;
        pixel_data[199][69] = 9;
        pixel_data[199][70] = 8;
        pixel_data[199][71] = 8;
        pixel_data[199][72] = 8;
        pixel_data[199][73] = 7;
        pixel_data[199][74] = 7;
        pixel_data[199][75] = 8;
        pixel_data[199][76] = 8;
        pixel_data[199][77] = 9;
        pixel_data[199][78] = 9;
        pixel_data[199][79] = 11;
        pixel_data[199][80] = 11;
        pixel_data[199][81] = 11;
        pixel_data[199][82] = 11;
        pixel_data[199][83] = 11;
        pixel_data[199][84] = 0;
        pixel_data[199][85] = 0;
        pixel_data[199][86] = 0;
        pixel_data[199][87] = 0;
        pixel_data[199][88] = 0;
        pixel_data[199][89] = 0;
        pixel_data[199][90] = 0;
        pixel_data[199][91] = 0;
        pixel_data[199][92] = 0;
        pixel_data[199][93] = 0;
        pixel_data[199][94] = 0;
        pixel_data[199][95] = 0;
        pixel_data[199][96] = 0;
        pixel_data[199][97] = 0;
        pixel_data[199][98] = 0;
        pixel_data[199][99] = 0;
        pixel_data[199][100] = 0;
        pixel_data[199][101] = 0;
        pixel_data[199][102] = 0;
        pixel_data[199][103] = 0;
        pixel_data[199][104] = 0;
        pixel_data[199][105] = 0;
        pixel_data[199][106] = 0;
        pixel_data[199][107] = 0;
        pixel_data[199][108] = 0;
        pixel_data[199][109] = 0;
        pixel_data[199][110] = 0;
        pixel_data[199][111] = 0;
        pixel_data[199][112] = 0;
        pixel_data[199][113] = 0;
        pixel_data[199][114] = 0;
        pixel_data[199][115] = 0;
        pixel_data[199][116] = 0;
        pixel_data[199][117] = 0;
        pixel_data[199][118] = 0;
        pixel_data[199][119] = 0;
        pixel_data[199][120] = 0;
        pixel_data[199][121] = 0;
        pixel_data[199][122] = 0;
        pixel_data[199][123] = 0;
        pixel_data[199][124] = 0;
        pixel_data[199][125] = 0;
        pixel_data[199][126] = 0;
        pixel_data[199][127] = 0;
        pixel_data[199][128] = 0;
        pixel_data[199][129] = 0;
        pixel_data[199][130] = 0;
        pixel_data[199][131] = 0;
        pixel_data[199][132] = 0;
        pixel_data[199][133] = 0;
        pixel_data[199][134] = 0;
        pixel_data[199][135] = 0;
        pixel_data[199][136] = 0;
        pixel_data[199][137] = 0;
        pixel_data[199][138] = 0;
        pixel_data[199][139] = 0;
        pixel_data[199][140] = 0;
        pixel_data[199][141] = 0;
        pixel_data[199][142] = 0;
        pixel_data[199][143] = 0;
        pixel_data[199][144] = 0;
        pixel_data[199][145] = 0;
        pixel_data[199][146] = 0;
        pixel_data[199][147] = 0;
        pixel_data[199][148] = 0;
        pixel_data[199][149] = 0;
        pixel_data[199][150] = 0;
        pixel_data[199][151] = 0;
        pixel_data[199][152] = 0;
        pixel_data[199][153] = 0;
        pixel_data[199][154] = 0;
        pixel_data[199][155] = 0;
        pixel_data[199][156] = 0;
        pixel_data[199][157] = 0;
        pixel_data[199][158] = 0;
        pixel_data[199][159] = 0;
        pixel_data[199][160] = 0;
        pixel_data[199][161] = 0;
        pixel_data[199][162] = 0;
        pixel_data[199][163] = 0;
        pixel_data[199][164] = 0;
        pixel_data[199][165] = 0;
        pixel_data[199][166] = 0;
        pixel_data[199][167] = 0;
        pixel_data[199][168] = 0;
        pixel_data[199][169] = 0;
        pixel_data[199][170] = 0;
        pixel_data[199][171] = 0;
        pixel_data[199][172] = 0;
        pixel_data[199][173] = 0;
        pixel_data[199][174] = 0;
        pixel_data[199][175] = 0;
        pixel_data[199][176] = 0;
        pixel_data[199][177] = 0;
        pixel_data[199][178] = 0;
        pixel_data[199][179] = 0;
        pixel_data[199][180] = 0;
        pixel_data[199][181] = 0;
        pixel_data[199][182] = 0;
        pixel_data[199][183] = 0;
        pixel_data[199][184] = 0;
        pixel_data[199][185] = 0;
        pixel_data[199][186] = 0;
        pixel_data[199][187] = 0;
        pixel_data[199][188] = 0;
        pixel_data[199][189] = 0;
        pixel_data[199][190] = 0;
        pixel_data[199][191] = 0;
        pixel_data[199][192] = 0;
        pixel_data[199][193] = 0;
        pixel_data[199][194] = 0;
        pixel_data[199][195] = 0;
        pixel_data[199][196] = 0;
        pixel_data[199][197] = 0;
        pixel_data[199][198] = 0;
        pixel_data[199][199] = 0; // y=199
    end
endmodule
