package SramPkg;
   localparam int MAP_X = 1023; // Maximum X coordinate
   localparam int MAP_Y = 767;  // Maximum Y coordinate
   localparam int PLAYER_X = 512; // Player's initial X coordinate
   localparam int PLAYER_Y = 384; // Player's initial Y coordinate
   localparam int SQUAT_PLAYER_Y = 512; // Player's initial Y coordinate
   localparam int BULLET_X = 512; // Bullet's initial X coordinate
   localparam int BULLET_Y = 384; // Bullet's initial Y coordinate
endpackage
