module player2_shield_palette(output reg [23:0] color_map [0:15]);
    initial begin
        color_map[0] = 24'h000000; // Transparent
        color_map[1] = 24'hfefe00;
        color_map[2] = 24'h90f64f;
        color_map[3] = 24'h7de13d;
        color_map[4] = 24'ha5b13c;
        color_map[5] = 24'hff7f00;
        color_map[6] = 24'hc48239;
        color_map[7] = 24'hc67d37;
        color_map[8] = 24'hd1625d;
        color_map[9] = 24'he64e7e;
        color_map[10] = 24'hb46e3a;
        color_map[11] = 24'he94d35;
        color_map[12] = 24'hed412d;
        color_map[13] = 24'hf12a0f;
        color_map[14] = 24'h814921;
        color_map[15] = 24'hfe0000;
    end
endmodule

module player2_shield_lut(output reg [3:0] pixel_data [0:49][0:49]);
    initial begin
        pixel_data[0][0] = 0;
        pixel_data[0][1] = 0;
        pixel_data[0][2] = 0;
        pixel_data[0][3] = 0;
        pixel_data[0][4] = 0;
        pixel_data[0][5] = 0;
        pixel_data[0][6] = 0;
        pixel_data[0][7] = 0;
        pixel_data[0][8] = 0;
        pixel_data[0][9] = 0;
        pixel_data[0][10] = 0;
        pixel_data[0][11] = 0;
        pixel_data[0][12] = 0;
        pixel_data[0][13] = 0;
        pixel_data[0][14] = 0;
        pixel_data[0][15] = 1;
        pixel_data[0][16] = 9;
        pixel_data[0][17] = 0;
        pixel_data[0][18] = 0;
        pixel_data[0][19] = 0;
        pixel_data[0][20] = 0;
        pixel_data[0][21] = 1;
        pixel_data[0][22] = 11;
        pixel_data[0][23] = 11;
        pixel_data[0][24] = 1;
        pixel_data[0][25] = 1;
        pixel_data[0][26] = 1;
        pixel_data[0][27] = 11;
        pixel_data[0][28] = 7;
        pixel_data[0][29] = 4;
        pixel_data[0][30] = 15;
        pixel_data[0][31] = 13;
        pixel_data[0][32] = 14;
        pixel_data[0][33] = 14;
        pixel_data[0][34] = 0;
        pixel_data[0][35] = 0;
        pixel_data[0][36] = 0;
        pixel_data[0][37] = 0;
        pixel_data[0][38] = 3;
        pixel_data[0][39] = 15;
        pixel_data[0][40] = 12;
        pixel_data[0][41] = 0;
        pixel_data[0][42] = 0;
        pixel_data[0][43] = 0;
        pixel_data[0][44] = 0;
        pixel_data[0][45] = 0;
        pixel_data[0][46] = 0;
        pixel_data[0][47] = 0;
        pixel_data[0][48] = 0;
        pixel_data[0][49] = 0; // y=0
        pixel_data[1][0] = 0;
        pixel_data[1][1] = 0;
        pixel_data[1][2] = 0;
        pixel_data[1][3] = 0;
        pixel_data[1][4] = 0;
        pixel_data[1][5] = 0;
        pixel_data[1][6] = 0;
        pixel_data[1][7] = 0;
        pixel_data[1][8] = 0;
        pixel_data[1][9] = 0;
        pixel_data[1][10] = 0;
        pixel_data[1][11] = 0;
        pixel_data[1][12] = 0;
        pixel_data[1][13] = 1;
        pixel_data[1][14] = 5;
        pixel_data[1][15] = 0;
        pixel_data[1][16] = 0;
        pixel_data[1][17] = 0;
        pixel_data[1][18] = 11;
        pixel_data[1][19] = 11;
        pixel_data[1][20] = 11;
        pixel_data[1][21] = 11;
        pixel_data[1][22] = 1;
        pixel_data[1][23] = 1;
        pixel_data[1][24] = 11;
        pixel_data[1][25] = 7;
        pixel_data[1][26] = 7;
        pixel_data[1][27] = 7;
        pixel_data[1][28] = 6;
        pixel_data[1][29] = 6;
        pixel_data[1][30] = 6;
        pixel_data[1][31] = 6;
        pixel_data[1][32] = 4;
        pixel_data[1][33] = 15;
        pixel_data[1][34] = 3;
        pixel_data[1][35] = 13;
        pixel_data[1][36] = 13;
        pixel_data[1][37] = 15;
        pixel_data[1][38] = 0;
        pixel_data[1][39] = 0;
        pixel_data[1][40] = 0;
        pixel_data[1][41] = 3;
        pixel_data[1][42] = 14;
        pixel_data[1][43] = 14;
        pixel_data[1][44] = 12;
        pixel_data[1][45] = 0;
        pixel_data[1][46] = 0;
        pixel_data[1][47] = 0;
        pixel_data[1][48] = 0;
        pixel_data[1][49] = 0; // y=1
        pixel_data[2][0] = 0;
        pixel_data[2][1] = 0;
        pixel_data[2][2] = 0;
        pixel_data[2][3] = 0;
        pixel_data[2][4] = 0;
        pixel_data[2][5] = 0;
        pixel_data[2][6] = 0;
        pixel_data[2][7] = 0;
        pixel_data[2][8] = 0;
        pixel_data[2][9] = 0;
        pixel_data[2][10] = 0;
        pixel_data[2][11] = 0;
        pixel_data[2][12] = 5;
        pixel_data[2][13] = 0;
        pixel_data[2][14] = 0;
        pixel_data[2][15] = 11;
        pixel_data[2][16] = 11;
        pixel_data[2][17] = 11;
        pixel_data[2][18] = 11;
        pixel_data[2][19] = 11;
        pixel_data[2][20] = 11;
        pixel_data[2][21] = 1;
        pixel_data[2][22] = 11;
        pixel_data[2][23] = 7;
        pixel_data[2][24] = 6;
        pixel_data[2][25] = 6;
        pixel_data[2][26] = 6;
        pixel_data[2][27] = 6;
        pixel_data[2][28] = 6;
        pixel_data[2][29] = 6;
        pixel_data[2][30] = 7;
        pixel_data[2][31] = 7;
        pixel_data[2][32] = 7;
        pixel_data[2][33] = 6;
        pixel_data[2][34] = 6;
        pixel_data[2][35] = 15;
        pixel_data[2][36] = 15;
        pixel_data[2][37] = 13;
        pixel_data[2][38] = 13;
        pixel_data[2][39] = 3;
        pixel_data[2][40] = 13;
        pixel_data[2][41] = 0;
        pixel_data[2][42] = 0;
        pixel_data[2][43] = 0;
        pixel_data[2][44] = 0;
        pixel_data[2][45] = 14;
        pixel_data[2][46] = 0;
        pixel_data[2][47] = 0;
        pixel_data[2][48] = 0;
        pixel_data[2][49] = 0; // y=2
        pixel_data[3][0] = 0;
        pixel_data[3][1] = 0;
        pixel_data[3][2] = 0;
        pixel_data[3][3] = 0;
        pixel_data[3][4] = 0;
        pixel_data[3][5] = 0;
        pixel_data[3][6] = 0;
        pixel_data[3][7] = 0;
        pixel_data[3][8] = 0;
        pixel_data[3][9] = 0;
        pixel_data[3][10] = 1;
        pixel_data[3][11] = 7;
        pixel_data[3][12] = 0;
        pixel_data[3][13] = 1;
        pixel_data[3][14] = 11;
        pixel_data[3][15] = 11;
        pixel_data[3][16] = 11;
        pixel_data[3][17] = 11;
        pixel_data[3][18] = 11;
        pixel_data[3][19] = 1;
        pixel_data[3][20] = 11;
        pixel_data[3][21] = 7;
        pixel_data[3][22] = 6;
        pixel_data[3][23] = 6;
        pixel_data[3][24] = 6;
        pixel_data[3][25] = 6;
        pixel_data[3][26] = 6;
        pixel_data[3][27] = 6;
        pixel_data[3][28] = 6;
        pixel_data[3][29] = 6;
        pixel_data[3][30] = 6;
        pixel_data[3][31] = 6;
        pixel_data[3][32] = 6;
        pixel_data[3][33] = 6;
        pixel_data[3][34] = 7;
        pixel_data[3][35] = 7;
        pixel_data[3][36] = 6;
        pixel_data[3][37] = 4;
        pixel_data[3][38] = 13;
        pixel_data[3][39] = 13;
        pixel_data[3][40] = 13;
        pixel_data[3][41] = 13;
        pixel_data[3][42] = 13;
        pixel_data[3][43] = 13;
        pixel_data[3][44] = 13;
        pixel_data[3][45] = 0;
        pixel_data[3][46] = 0;
        pixel_data[3][47] = 0;
        pixel_data[3][48] = 0;
        pixel_data[3][49] = 0; // y=3
        pixel_data[4][0] = 0;
        pixel_data[4][1] = 0;
        pixel_data[4][2] = 0;
        pixel_data[4][3] = 0;
        pixel_data[4][4] = 0;
        pixel_data[4][5] = 0;
        pixel_data[4][6] = 0;
        pixel_data[4][7] = 0;
        pixel_data[4][8] = 0;
        pixel_data[4][9] = 5;
        pixel_data[4][10] = 0;
        pixel_data[4][11] = 0;
        pixel_data[4][12] = 11;
        pixel_data[4][13] = 11;
        pixel_data[4][14] = 11;
        pixel_data[4][15] = 11;
        pixel_data[4][16] = 11;
        pixel_data[4][17] = 11;
        pixel_data[4][18] = 1;
        pixel_data[4][19] = 11;
        pixel_data[4][20] = 7;
        pixel_data[4][21] = 6;
        pixel_data[4][22] = 6;
        pixel_data[4][23] = 6;
        pixel_data[4][24] = 6;
        pixel_data[4][25] = 6;
        pixel_data[4][26] = 6;
        pixel_data[4][27] = 6;
        pixel_data[4][28] = 6;
        pixel_data[4][29] = 6;
        pixel_data[4][30] = 6;
        pixel_data[4][31] = 6;
        pixel_data[4][32] = 6;
        pixel_data[4][33] = 6;
        pixel_data[4][34] = 6;
        pixel_data[4][35] = 6;
        pixel_data[4][36] = 6;
        pixel_data[4][37] = 7;
        pixel_data[4][38] = 6;
        pixel_data[4][39] = 15;
        pixel_data[4][40] = 13;
        pixel_data[4][41] = 13;
        pixel_data[4][42] = 13;
        pixel_data[4][43] = 13;
        pixel_data[4][44] = 13;
        pixel_data[4][45] = 13;
        pixel_data[4][46] = 0;
        pixel_data[4][47] = 14;
        pixel_data[4][48] = 0;
        pixel_data[4][49] = 0; // y=4
        pixel_data[5][0] = 0;
        pixel_data[5][1] = 0;
        pixel_data[5][2] = 0;
        pixel_data[5][3] = 0;
        pixel_data[5][4] = 0;
        pixel_data[5][5] = 0;
        pixel_data[5][6] = 0;
        pixel_data[5][7] = 0;
        pixel_data[5][8] = 5;
        pixel_data[5][9] = 0;
        pixel_data[5][10] = 11;
        pixel_data[5][11] = 1;
        pixel_data[5][12] = 1;
        pixel_data[5][13] = 1;
        pixel_data[5][14] = 1;
        pixel_data[5][15] = 11;
        pixel_data[5][16] = 11;
        pixel_data[5][17] = 1;
        pixel_data[5][18] = 7;
        pixel_data[5][19] = 6;
        pixel_data[5][20] = 6;
        pixel_data[5][21] = 6;
        pixel_data[5][22] = 6;
        pixel_data[5][23] = 6;
        pixel_data[5][24] = 6;
        pixel_data[5][25] = 6;
        pixel_data[5][26] = 6;
        pixel_data[5][27] = 6;
        pixel_data[5][28] = 6;
        pixel_data[5][29] = 6;
        pixel_data[5][30] = 6;
        pixel_data[5][31] = 6;
        pixel_data[5][32] = 6;
        pixel_data[5][33] = 6;
        pixel_data[5][34] = 6;
        pixel_data[5][35] = 6;
        pixel_data[5][36] = 6;
        pixel_data[5][37] = 6;
        pixel_data[5][38] = 7;
        pixel_data[5][39] = 7;
        pixel_data[5][40] = 4;
        pixel_data[5][41] = 3;
        pixel_data[5][42] = 13;
        pixel_data[5][43] = 13;
        pixel_data[5][44] = 13;
        pixel_data[5][45] = 13;
        pixel_data[5][46] = 0;
        pixel_data[5][47] = 14;
        pixel_data[5][48] = 0;
        pixel_data[5][49] = 0; // y=5
        pixel_data[6][0] = 0;
        pixel_data[6][1] = 0;
        pixel_data[6][2] = 0;
        pixel_data[6][3] = 0;
        pixel_data[6][4] = 0;
        pixel_data[6][5] = 0;
        pixel_data[6][6] = 0;
        pixel_data[6][7] = 5;
        pixel_data[6][8] = 0;
        pixel_data[6][9] = 11;
        pixel_data[6][10] = 1;
        pixel_data[6][11] = 1;
        pixel_data[6][12] = 1;
        pixel_data[6][13] = 1;
        pixel_data[6][14] = 1;
        pixel_data[6][15] = 11;
        pixel_data[6][16] = 11;
        pixel_data[6][17] = 7;
        pixel_data[6][18] = 6;
        pixel_data[6][19] = 6;
        pixel_data[6][20] = 6;
        pixel_data[6][21] = 6;
        pixel_data[6][22] = 6;
        pixel_data[6][23] = 6;
        pixel_data[6][24] = 6;
        pixel_data[6][25] = 6;
        pixel_data[6][26] = 6;
        pixel_data[6][27] = 6;
        pixel_data[6][28] = 6;
        pixel_data[6][29] = 6;
        pixel_data[6][30] = 6;
        pixel_data[6][31] = 6;
        pixel_data[6][32] = 6;
        pixel_data[6][33] = 6;
        pixel_data[6][34] = 6;
        pixel_data[6][35] = 6;
        pixel_data[6][36] = 6;
        pixel_data[6][37] = 6;
        pixel_data[6][38] = 6;
        pixel_data[6][39] = 7;
        pixel_data[6][40] = 11;
        pixel_data[6][41] = 11;
        pixel_data[6][42] = 11;
        pixel_data[6][43] = 13;
        pixel_data[6][44] = 12;
        pixel_data[6][45] = 13;
        pixel_data[6][46] = 0;
        pixel_data[6][47] = 14;
        pixel_data[6][48] = 0;
        pixel_data[6][49] = 0; // y=6
        pixel_data[7][0] = 0;
        pixel_data[7][1] = 0;
        pixel_data[7][2] = 0;
        pixel_data[7][3] = 0;
        pixel_data[7][4] = 0;
        pixel_data[7][5] = 0;
        pixel_data[7][6] = 14;
        pixel_data[7][7] = 0;
        pixel_data[7][8] = 11;
        pixel_data[7][9] = 1;
        pixel_data[7][10] = 1;
        pixel_data[7][11] = 1;
        pixel_data[7][12] = 1;
        pixel_data[7][13] = 1;
        pixel_data[7][14] = 1;
        pixel_data[7][15] = 11;
        pixel_data[7][16] = 7;
        pixel_data[7][17] = 6;
        pixel_data[7][18] = 6;
        pixel_data[7][19] = 6;
        pixel_data[7][20] = 6;
        pixel_data[7][21] = 6;
        pixel_data[7][22] = 6;
        pixel_data[7][23] = 6;
        pixel_data[7][24] = 6;
        pixel_data[7][25] = 6;
        pixel_data[7][26] = 6;
        pixel_data[7][27] = 6;
        pixel_data[7][28] = 6;
        pixel_data[7][29] = 6;
        pixel_data[7][30] = 6;
        pixel_data[7][31] = 6;
        pixel_data[7][32] = 6;
        pixel_data[7][33] = 6;
        pixel_data[7][34] = 6;
        pixel_data[7][35] = 6;
        pixel_data[7][36] = 6;
        pixel_data[7][37] = 6;
        pixel_data[7][38] = 6;
        pixel_data[7][39] = 11;
        pixel_data[7][40] = 1;
        pixel_data[7][41] = 11;
        pixel_data[7][42] = 1;
        pixel_data[7][43] = 4;
        pixel_data[7][44] = 13;
        pixel_data[7][45] = 15;
        pixel_data[7][46] = 0;
        pixel_data[7][47] = 12;
        pixel_data[7][48] = 0;
        pixel_data[7][49] = 0; // y=7
        pixel_data[8][0] = 0;
        pixel_data[8][1] = 0;
        pixel_data[8][2] = 0;
        pixel_data[8][3] = 0;
        pixel_data[8][4] = 0;
        pixel_data[8][5] = 5;
        pixel_data[8][6] = 0;
        pixel_data[8][7] = 11;
        pixel_data[8][8] = 11;
        pixel_data[8][9] = 1;
        pixel_data[8][10] = 1;
        pixel_data[8][11] = 1;
        pixel_data[8][12] = 1;
        pixel_data[8][13] = 1;
        pixel_data[8][14] = 11;
        pixel_data[8][15] = 7;
        pixel_data[8][16] = 6;
        pixel_data[8][17] = 6;
        pixel_data[8][18] = 6;
        pixel_data[8][19] = 6;
        pixel_data[8][20] = 6;
        pixel_data[8][21] = 6;
        pixel_data[8][22] = 6;
        pixel_data[8][23] = 6;
        pixel_data[8][24] = 6;
        pixel_data[8][25] = 6;
        pixel_data[8][26] = 6;
        pixel_data[8][27] = 6;
        pixel_data[8][28] = 6;
        pixel_data[8][29] = 6;
        pixel_data[8][30] = 6;
        pixel_data[8][31] = 6;
        pixel_data[8][32] = 6;
        pixel_data[8][33] = 6;
        pixel_data[8][34] = 6;
        pixel_data[8][35] = 6;
        pixel_data[8][36] = 6;
        pixel_data[8][37] = 6;
        pixel_data[8][38] = 7;
        pixel_data[8][39] = 1;
        pixel_data[8][40] = 11;
        pixel_data[8][41] = 11;
        pixel_data[8][42] = 11;
        pixel_data[8][43] = 1;
        pixel_data[8][44] = 0;
        pixel_data[8][45] = 0;
        pixel_data[8][46] = 1;
        pixel_data[8][47] = 0;
        pixel_data[8][48] = 0;
        pixel_data[8][49] = 0; // y=8
        pixel_data[9][0] = 0;
        pixel_data[9][1] = 0;
        pixel_data[9][2] = 0;
        pixel_data[9][3] = 0;
        pixel_data[9][4] = 5;
        pixel_data[9][5] = 0;
        pixel_data[9][6] = 11;
        pixel_data[9][7] = 11;
        pixel_data[9][8] = 11;
        pixel_data[9][9] = 1;
        pixel_data[9][10] = 1;
        pixel_data[9][11] = 1;
        pixel_data[9][12] = 1;
        pixel_data[9][13] = 1;
        pixel_data[9][14] = 7;
        pixel_data[9][15] = 6;
        pixel_data[9][16] = 6;
        pixel_data[9][17] = 6;
        pixel_data[9][18] = 6;
        pixel_data[9][19] = 6;
        pixel_data[9][20] = 6;
        pixel_data[9][21] = 6;
        pixel_data[9][22] = 6;
        pixel_data[9][23] = 6;
        pixel_data[9][24] = 6;
        pixel_data[9][25] = 6;
        pixel_data[9][26] = 6;
        pixel_data[9][27] = 6;
        pixel_data[9][28] = 6;
        pixel_data[9][29] = 6;
        pixel_data[9][30] = 6;
        pixel_data[9][31] = 6;
        pixel_data[9][32] = 6;
        pixel_data[9][33] = 6;
        pixel_data[9][34] = 6;
        pixel_data[9][35] = 6;
        pixel_data[9][36] = 6;
        pixel_data[9][37] = 7;
        pixel_data[9][38] = 11;
        pixel_data[9][39] = 11;
        pixel_data[9][40] = 11;
        pixel_data[9][41] = 11;
        pixel_data[9][42] = 11;
        pixel_data[9][43] = 11;
        pixel_data[9][44] = 11;
        pixel_data[9][45] = 9;
        pixel_data[9][46] = 5;
        pixel_data[9][47] = 0;
        pixel_data[9][48] = 0;
        pixel_data[9][49] = 0; // y=9
        pixel_data[10][0] = 0;
        pixel_data[10][1] = 0;
        pixel_data[10][2] = 0;
        pixel_data[10][3] = 1;
        pixel_data[10][4] = 0;
        pixel_data[10][5] = 11;
        pixel_data[10][6] = 11;
        pixel_data[10][7] = 1;
        pixel_data[10][8] = 1;
        pixel_data[10][9] = 11;
        pixel_data[10][10] = 1;
        pixel_data[10][11] = 11;
        pixel_data[10][12] = 1;
        pixel_data[10][13] = 11;
        pixel_data[10][14] = 6;
        pixel_data[10][15] = 6;
        pixel_data[10][16] = 6;
        pixel_data[10][17] = 6;
        pixel_data[10][18] = 6;
        pixel_data[10][19] = 6;
        pixel_data[10][20] = 6;
        pixel_data[10][21] = 6;
        pixel_data[10][22] = 6;
        pixel_data[10][23] = 6;
        pixel_data[10][24] = 6;
        pixel_data[10][25] = 6;
        pixel_data[10][26] = 6;
        pixel_data[10][27] = 6;
        pixel_data[10][28] = 6;
        pixel_data[10][29] = 6;
        pixel_data[10][30] = 6;
        pixel_data[10][31] = 6;
        pixel_data[10][32] = 6;
        pixel_data[10][33] = 6;
        pixel_data[10][34] = 6;
        pixel_data[10][35] = 6;
        pixel_data[10][36] = 6;
        pixel_data[10][37] = 7;
        pixel_data[10][38] = 1;
        pixel_data[10][39] = 11;
        pixel_data[10][40] = 11;
        pixel_data[10][41] = 11;
        pixel_data[10][42] = 11;
        pixel_data[10][43] = 11;
        pixel_data[10][44] = 11;
        pixel_data[10][45] = 11;
        pixel_data[10][46] = 0;
        pixel_data[10][47] = 5;
        pixel_data[10][48] = 0;
        pixel_data[10][49] = 0; // y=10
        pixel_data[11][0] = 0;
        pixel_data[11][1] = 0;
        pixel_data[11][2] = 1;
        pixel_data[11][3] = 3;
        pixel_data[11][4] = 11;
        pixel_data[11][5] = 11;
        pixel_data[11][6] = 1;
        pixel_data[11][7] = 1;
        pixel_data[11][8] = 1;
        pixel_data[11][9] = 1;
        pixel_data[11][10] = 11;
        pixel_data[11][11] = 1;
        pixel_data[11][12] = 11;
        pixel_data[11][13] = 7;
        pixel_data[11][14] = 6;
        pixel_data[11][15] = 6;
        pixel_data[11][16] = 6;
        pixel_data[11][17] = 6;
        pixel_data[11][18] = 6;
        pixel_data[11][19] = 6;
        pixel_data[11][20] = 6;
        pixel_data[11][21] = 6;
        pixel_data[11][22] = 6;
        pixel_data[11][23] = 6;
        pixel_data[11][24] = 6;
        pixel_data[11][25] = 6;
        pixel_data[11][26] = 6;
        pixel_data[11][27] = 6;
        pixel_data[11][28] = 6;
        pixel_data[11][29] = 6;
        pixel_data[11][30] = 6;
        pixel_data[11][31] = 6;
        pixel_data[11][32] = 6;
        pixel_data[11][33] = 6;
        pixel_data[11][34] = 6;
        pixel_data[11][35] = 6;
        pixel_data[11][36] = 6;
        pixel_data[11][37] = 11;
        pixel_data[11][38] = 1;
        pixel_data[11][39] = 11;
        pixel_data[11][40] = 11;
        pixel_data[11][41] = 11;
        pixel_data[11][42] = 11;
        pixel_data[11][43] = 11;
        pixel_data[11][44] = 11;
        pixel_data[11][45] = 11;
        pixel_data[11][46] = 11;
        pixel_data[11][47] = 0;
        pixel_data[11][48] = 1;
        pixel_data[11][49] = 0; // y=11
        pixel_data[12][0] = 0;
        pixel_data[12][1] = 0;
        pixel_data[12][2] = 5;
        pixel_data[12][3] = 0;
        pixel_data[12][4] = 11;
        pixel_data[12][5] = 1;
        pixel_data[12][6] = 1;
        pixel_data[12][7] = 1;
        pixel_data[12][8] = 1;
        pixel_data[12][9] = 1;
        pixel_data[12][10] = 11;
        pixel_data[12][11] = 11;
        pixel_data[12][12] = 7;
        pixel_data[12][13] = 6;
        pixel_data[12][14] = 6;
        pixel_data[12][15] = 6;
        pixel_data[12][16] = 6;
        pixel_data[12][17] = 6;
        pixel_data[12][18] = 6;
        pixel_data[12][19] = 6;
        pixel_data[12][20] = 6;
        pixel_data[12][21] = 6;
        pixel_data[12][22] = 6;
        pixel_data[12][23] = 6;
        pixel_data[12][24] = 6;
        pixel_data[12][25] = 6;
        pixel_data[12][26] = 6;
        pixel_data[12][27] = 6;
        pixel_data[12][28] = 6;
        pixel_data[12][29] = 6;
        pixel_data[12][30] = 6;
        pixel_data[12][31] = 6;
        pixel_data[12][32] = 6;
        pixel_data[12][33] = 6;
        pixel_data[12][34] = 6;
        pixel_data[12][35] = 6;
        pixel_data[12][36] = 6;
        pixel_data[12][37] = 11;
        pixel_data[12][38] = 11;
        pixel_data[12][39] = 11;
        pixel_data[12][40] = 11;
        pixel_data[12][41] = 11;
        pixel_data[12][42] = 11;
        pixel_data[12][43] = 11;
        pixel_data[12][44] = 11;
        pixel_data[12][45] = 11;
        pixel_data[12][46] = 11;
        pixel_data[12][47] = 0;
        pixel_data[12][48] = 12;
        pixel_data[12][49] = 0; // y=12
        pixel_data[13][0] = 0;
        pixel_data[13][1] = 1;
        pixel_data[13][2] = 0;
        pixel_data[13][3] = 11;
        pixel_data[13][4] = 1;
        pixel_data[13][5] = 1;
        pixel_data[13][6] = 1;
        pixel_data[13][7] = 1;
        pixel_data[13][8] = 1;
        pixel_data[13][9] = 11;
        pixel_data[13][10] = 1;
        pixel_data[13][11] = 7;
        pixel_data[13][12] = 6;
        pixel_data[13][13] = 6;
        pixel_data[13][14] = 6;
        pixel_data[13][15] = 6;
        pixel_data[13][16] = 6;
        pixel_data[13][17] = 6;
        pixel_data[13][18] = 6;
        pixel_data[13][19] = 6;
        pixel_data[13][20] = 6;
        pixel_data[13][21] = 6;
        pixel_data[13][22] = 6;
        pixel_data[13][23] = 6;
        pixel_data[13][24] = 6;
        pixel_data[13][25] = 6;
        pixel_data[13][26] = 6;
        pixel_data[13][27] = 6;
        pixel_data[13][28] = 6;
        pixel_data[13][29] = 6;
        pixel_data[13][30] = 6;
        pixel_data[13][31] = 6;
        pixel_data[13][32] = 6;
        pixel_data[13][33] = 6;
        pixel_data[13][34] = 6;
        pixel_data[13][35] = 6;
        pixel_data[13][36] = 6;
        pixel_data[13][37] = 11;
        pixel_data[13][38] = 11;
        pixel_data[13][39] = 11;
        pixel_data[13][40] = 11;
        pixel_data[13][41] = 11;
        pixel_data[13][42] = 11;
        pixel_data[13][43] = 11;
        pixel_data[13][44] = 11;
        pixel_data[13][45] = 11;
        pixel_data[13][46] = 11;
        pixel_data[13][47] = 11;
        pixel_data[13][48] = 0;
        pixel_data[13][49] = 5; // y=13
        pixel_data[14][0] = 0;
        pixel_data[14][1] = 1;
        pixel_data[14][2] = 0;
        pixel_data[14][3] = 1;
        pixel_data[14][4] = 1;
        pixel_data[14][5] = 1;
        pixel_data[14][6] = 1;
        pixel_data[14][7] = 1;
        pixel_data[14][8] = 1;
        pixel_data[14][9] = 1;
        pixel_data[14][10] = 11;
        pixel_data[14][11] = 6;
        pixel_data[14][12] = 6;
        pixel_data[14][13] = 6;
        pixel_data[14][14] = 6;
        pixel_data[14][15] = 6;
        pixel_data[14][16] = 6;
        pixel_data[14][17] = 6;
        pixel_data[14][18] = 6;
        pixel_data[14][19] = 6;
        pixel_data[14][20] = 6;
        pixel_data[14][21] = 6;
        pixel_data[14][22] = 6;
        pixel_data[14][23] = 6;
        pixel_data[14][24] = 6;
        pixel_data[14][25] = 6;
        pixel_data[14][26] = 6;
        pixel_data[14][27] = 6;
        pixel_data[14][28] = 6;
        pixel_data[14][29] = 6;
        pixel_data[14][30] = 6;
        pixel_data[14][31] = 6;
        pixel_data[14][32] = 6;
        pixel_data[14][33] = 6;
        pixel_data[14][34] = 6;
        pixel_data[14][35] = 6;
        pixel_data[14][36] = 6;
        pixel_data[14][37] = 11;
        pixel_data[14][38] = 1;
        pixel_data[14][39] = 11;
        pixel_data[14][40] = 11;
        pixel_data[14][41] = 11;
        pixel_data[14][42] = 11;
        pixel_data[14][43] = 11;
        pixel_data[14][44] = 11;
        pixel_data[14][45] = 11;
        pixel_data[14][46] = 11;
        pixel_data[14][47] = 11;
        pixel_data[14][48] = 0;
        pixel_data[14][49] = 14; // y=14
        pixel_data[15][0] = 1;
        pixel_data[15][1] = 0;
        pixel_data[15][2] = 1;
        pixel_data[15][3] = 1;
        pixel_data[15][4] = 1;
        pixel_data[15][5] = 1;
        pixel_data[15][6] = 1;
        pixel_data[15][7] = 1;
        pixel_data[15][8] = 11;
        pixel_data[15][9] = 1;
        pixel_data[15][10] = 7;
        pixel_data[15][11] = 6;
        pixel_data[15][12] = 6;
        pixel_data[15][13] = 6;
        pixel_data[15][14] = 6;
        pixel_data[15][15] = 6;
        pixel_data[15][16] = 6;
        pixel_data[15][17] = 6;
        pixel_data[15][18] = 6;
        pixel_data[15][19] = 6;
        pixel_data[15][20] = 6;
        pixel_data[15][21] = 6;
        pixel_data[15][22] = 6;
        pixel_data[15][23] = 6;
        pixel_data[15][24] = 6;
        pixel_data[15][25] = 6;
        pixel_data[15][26] = 7;
        pixel_data[15][27] = 7;
        pixel_data[15][28] = 6;
        pixel_data[15][29] = 6;
        pixel_data[15][30] = 6;
        pixel_data[15][31] = 6;
        pixel_data[15][32] = 6;
        pixel_data[15][33] = 6;
        pixel_data[15][34] = 6;
        pixel_data[15][35] = 6;
        pixel_data[15][36] = 6;
        pixel_data[15][37] = 11;
        pixel_data[15][38] = 1;
        pixel_data[15][39] = 11;
        pixel_data[15][40] = 11;
        pixel_data[15][41] = 11;
        pixel_data[15][42] = 11;
        pixel_data[15][43] = 11;
        pixel_data[15][44] = 11;
        pixel_data[15][45] = 11;
        pixel_data[15][46] = 11;
        pixel_data[15][47] = 11;
        pixel_data[15][48] = 1;
        pixel_data[15][49] = 0; // y=15
        pixel_data[16][0] = 1;
        pixel_data[16][1] = 0;
        pixel_data[16][2] = 1;
        pixel_data[16][3] = 1;
        pixel_data[16][4] = 1;
        pixel_data[16][5] = 1;
        pixel_data[16][6] = 1;
        pixel_data[16][7] = 11;
        pixel_data[16][8] = 1;
        pixel_data[16][9] = 11;
        pixel_data[16][10] = 6;
        pixel_data[16][11] = 7;
        pixel_data[16][12] = 7;
        pixel_data[16][13] = 6;
        pixel_data[16][14] = 6;
        pixel_data[16][15] = 8;
        pixel_data[16][16] = 8;
        pixel_data[16][17] = 8;
        pixel_data[16][18] = 6;
        pixel_data[16][19] = 6;
        pixel_data[16][20] = 6;
        pixel_data[16][21] = 6;
        pixel_data[16][22] = 6;
        pixel_data[16][23] = 6;
        pixel_data[16][24] = 6;
        pixel_data[16][25] = 8;
        pixel_data[16][26] = 9;
        pixel_data[16][27] = 9;
        pixel_data[16][28] = 9;
        pixel_data[16][29] = 8;
        pixel_data[16][30] = 6;
        pixel_data[16][31] = 6;
        pixel_data[16][32] = 6;
        pixel_data[16][33] = 6;
        pixel_data[16][34] = 6;
        pixel_data[16][35] = 6;
        pixel_data[16][36] = 6;
        pixel_data[16][37] = 7;
        pixel_data[16][38] = 1;
        pixel_data[16][39] = 11;
        pixel_data[16][40] = 11;
        pixel_data[16][41] = 11;
        pixel_data[16][42] = 11;
        pixel_data[16][43] = 11;
        pixel_data[16][44] = 11;
        pixel_data[16][45] = 11;
        pixel_data[16][46] = 11;
        pixel_data[16][47] = 11;
        pixel_data[16][48] = 11;
        pixel_data[16][49] = 0; // y=16
        pixel_data[17][0] = 0;
        pixel_data[17][1] = 1;
        pixel_data[17][2] = 1;
        pixel_data[17][3] = 1;
        pixel_data[17][4] = 1;
        pixel_data[17][5] = 1;
        pixel_data[17][6] = 1;
        pixel_data[17][7] = 11;
        pixel_data[17][8] = 11;
        pixel_data[17][9] = 7;
        pixel_data[17][10] = 6;
        pixel_data[17][11] = 7;
        pixel_data[17][12] = 7;
        pixel_data[17][13] = 7;
        pixel_data[17][14] = 9;
        pixel_data[17][15] = 9;
        pixel_data[17][16] = 9;
        pixel_data[17][17] = 1;
        pixel_data[17][18] = 8;
        pixel_data[17][19] = 6;
        pixel_data[17][20] = 6;
        pixel_data[17][21] = 6;
        pixel_data[17][22] = 6;
        pixel_data[17][23] = 6;
        pixel_data[17][24] = 7;
        pixel_data[17][25] = 9;
        pixel_data[17][26] = 9;
        pixel_data[17][27] = 9;
        pixel_data[17][28] = 9;
        pixel_data[17][29] = 9;
        pixel_data[17][30] = 8;
        pixel_data[17][31] = 6;
        pixel_data[17][32] = 6;
        pixel_data[17][33] = 6;
        pixel_data[17][34] = 6;
        pixel_data[17][35] = 6;
        pixel_data[17][36] = 6;
        pixel_data[17][37] = 7;
        pixel_data[17][38] = 11;
        pixel_data[17][39] = 11;
        pixel_data[17][40] = 11;
        pixel_data[17][41] = 11;
        pixel_data[17][42] = 11;
        pixel_data[17][43] = 11;
        pixel_data[17][44] = 11;
        pixel_data[17][45] = 11;
        pixel_data[17][46] = 11;
        pixel_data[17][47] = 11;
        pixel_data[17][48] = 11;
        pixel_data[17][49] = 0; // y=17
        pixel_data[18][0] = 0;
        pixel_data[18][1] = 1;
        pixel_data[18][2] = 1;
        pixel_data[18][3] = 1;
        pixel_data[18][4] = 1;
        pixel_data[18][5] = 1;
        pixel_data[18][6] = 11;
        pixel_data[18][7] = 1;
        pixel_data[18][8] = 7;
        pixel_data[18][9] = 6;
        pixel_data[18][10] = 7;
        pixel_data[18][11] = 10;
        pixel_data[18][12] = 10;
        pixel_data[18][13] = 9;
        pixel_data[18][14] = 9;
        pixel_data[18][15] = 9;
        pixel_data[18][16] = 9;
        pixel_data[18][17] = 9;
        pixel_data[18][18] = 9;
        pixel_data[18][19] = 6;
        pixel_data[18][20] = 6;
        pixel_data[18][21] = 6;
        pixel_data[18][22] = 6;
        pixel_data[18][23] = 6;
        pixel_data[18][24] = 8;
        pixel_data[18][25] = 9;
        pixel_data[18][26] = 9;
        pixel_data[18][27] = 9;
        pixel_data[18][28] = 9;
        pixel_data[18][29] = 9;
        pixel_data[18][30] = 9;
        pixel_data[18][31] = 8;
        pixel_data[18][32] = 6;
        pixel_data[18][33] = 6;
        pixel_data[18][34] = 6;
        pixel_data[18][35] = 6;
        pixel_data[18][36] = 6;
        pixel_data[18][37] = 6;
        pixel_data[18][38] = 11;
        pixel_data[18][39] = 1;
        pixel_data[18][40] = 11;
        pixel_data[18][41] = 11;
        pixel_data[18][42] = 11;
        pixel_data[18][43] = 11;
        pixel_data[18][44] = 11;
        pixel_data[18][45] = 11;
        pixel_data[18][46] = 11;
        pixel_data[18][47] = 11;
        pixel_data[18][48] = 11;
        pixel_data[18][49] = 11; // y=18
        pixel_data[19][0] = 0;
        pixel_data[19][1] = 1;
        pixel_data[19][2] = 1;
        pixel_data[19][3] = 1;
        pixel_data[19][4] = 1;
        pixel_data[19][5] = 1;
        pixel_data[19][6] = 11;
        pixel_data[19][7] = 11;
        pixel_data[19][8] = 6;
        pixel_data[19][9] = 7;
        pixel_data[19][10] = 7;
        pixel_data[19][11] = 10;
        pixel_data[19][12] = 8;
        pixel_data[19][13] = 9;
        pixel_data[19][14] = 9;
        pixel_data[19][15] = 9;
        pixel_data[19][16] = 9;
        pixel_data[19][17] = 9;
        pixel_data[19][18] = 9;
        pixel_data[19][19] = 6;
        pixel_data[19][20] = 6;
        pixel_data[19][21] = 6;
        pixel_data[19][22] = 6;
        pixel_data[19][23] = 6;
        pixel_data[19][24] = 8;
        pixel_data[19][25] = 9;
        pixel_data[19][26] = 9;
        pixel_data[19][27] = 9;
        pixel_data[19][28] = 9;
        pixel_data[19][29] = 9;
        pixel_data[19][30] = 9;
        pixel_data[19][31] = 9;
        pixel_data[19][32] = 8;
        pixel_data[19][33] = 6;
        pixel_data[19][34] = 10;
        pixel_data[19][35] = 7;
        pixel_data[19][36] = 6;
        pixel_data[19][37] = 6;
        pixel_data[19][38] = 7;
        pixel_data[19][39] = 1;
        pixel_data[19][40] = 11;
        pixel_data[19][41] = 11;
        pixel_data[19][42] = 11;
        pixel_data[19][43] = 11;
        pixel_data[19][44] = 11;
        pixel_data[19][45] = 11;
        pixel_data[19][46] = 11;
        pixel_data[19][47] = 11;
        pixel_data[19][48] = 11;
        pixel_data[19][49] = 11; // y=19
        pixel_data[20][0] = 1;
        pixel_data[20][1] = 1;
        pixel_data[20][2] = 1;
        pixel_data[20][3] = 1;
        pixel_data[20][4] = 1;
        pixel_data[20][5] = 1;
        pixel_data[20][6] = 1;
        pixel_data[20][7] = 7;
        pixel_data[20][8] = 6;
        pixel_data[20][9] = 7;
        pixel_data[20][10] = 10;
        pixel_data[20][11] = 10;
        pixel_data[20][12] = 9;
        pixel_data[20][13] = 9;
        pixel_data[20][14] = 9;
        pixel_data[20][15] = 9;
        pixel_data[20][16] = 9;
        pixel_data[20][17] = 9;
        pixel_data[20][18] = 8;
        pixel_data[20][19] = 6;
        pixel_data[20][20] = 6;
        pixel_data[20][21] = 6;
        pixel_data[20][22] = 6;
        pixel_data[20][23] = 6;
        pixel_data[20][24] = 9;
        pixel_data[20][25] = 9;
        pixel_data[20][26] = 9;
        pixel_data[20][27] = 9;
        pixel_data[20][28] = 9;
        pixel_data[20][29] = 9;
        pixel_data[20][30] = 9;
        pixel_data[20][31] = 9;
        pixel_data[20][32] = 9;
        pixel_data[20][33] = 7;
        pixel_data[20][34] = 10;
        pixel_data[20][35] = 10;
        pixel_data[20][36] = 6;
        pixel_data[20][37] = 6;
        pixel_data[20][38] = 6;
        pixel_data[20][39] = 11;
        pixel_data[20][40] = 11;
        pixel_data[20][41] = 11;
        pixel_data[20][42] = 11;
        pixel_data[20][43] = 11;
        pixel_data[20][44] = 11;
        pixel_data[20][45] = 11;
        pixel_data[20][46] = 11;
        pixel_data[20][47] = 11;
        pixel_data[20][48] = 11;
        pixel_data[20][49] = 11; // y=20
        pixel_data[21][0] = 1;
        pixel_data[21][1] = 1;
        pixel_data[21][2] = 1;
        pixel_data[21][3] = 1;
        pixel_data[21][4] = 1;
        pixel_data[21][5] = 1;
        pixel_data[21][6] = 11;
        pixel_data[21][7] = 7;
        pixel_data[21][8] = 7;
        pixel_data[21][9] = 7;
        pixel_data[21][10] = 10;
        pixel_data[21][11] = 8;
        pixel_data[21][12] = 9;
        pixel_data[21][13] = 9;
        pixel_data[21][14] = 9;
        pixel_data[21][15] = 9;
        pixel_data[21][16] = 9;
        pixel_data[21][17] = 9;
        pixel_data[21][18] = 8;
        pixel_data[21][19] = 6;
        pixel_data[21][20] = 6;
        pixel_data[21][21] = 6;
        pixel_data[21][22] = 6;
        pixel_data[21][23] = 6;
        pixel_data[21][24] = 9;
        pixel_data[21][25] = 9;
        pixel_data[21][26] = 9;
        pixel_data[21][27] = 9;
        pixel_data[21][28] = 9;
        pixel_data[21][29] = 9;
        pixel_data[21][30] = 9;
        pixel_data[21][31] = 9;
        pixel_data[21][32] = 9;
        pixel_data[21][33] = 8;
        pixel_data[21][34] = 10;
        pixel_data[21][35] = 10;
        pixel_data[21][36] = 6;
        pixel_data[21][37] = 6;
        pixel_data[21][38] = 6;
        pixel_data[21][39] = 7;
        pixel_data[21][40] = 1;
        pixel_data[21][41] = 11;
        pixel_data[21][42] = 11;
        pixel_data[21][43] = 11;
        pixel_data[21][44] = 11;
        pixel_data[21][45] = 11;
        pixel_data[21][46] = 11;
        pixel_data[21][47] = 11;
        pixel_data[21][48] = 11;
        pixel_data[21][49] = 1; // y=21
        pixel_data[22][0] = 1;
        pixel_data[22][1] = 1;
        pixel_data[22][2] = 1;
        pixel_data[22][3] = 1;
        pixel_data[22][4] = 1;
        pixel_data[22][5] = 1;
        pixel_data[22][6] = 7;
        pixel_data[22][7] = 7;
        pixel_data[22][8] = 7;
        pixel_data[22][9] = 10;
        pixel_data[22][10] = 10;
        pixel_data[22][11] = 9;
        pixel_data[22][12] = 9;
        pixel_data[22][13] = 9;
        pixel_data[22][14] = 9;
        pixel_data[22][15] = 9;
        pixel_data[22][16] = 9;
        pixel_data[22][17] = 8;
        pixel_data[22][18] = 7;
        pixel_data[22][19] = 6;
        pixel_data[22][20] = 6;
        pixel_data[22][21] = 6;
        pixel_data[22][22] = 6;
        pixel_data[22][23] = 6;
        pixel_data[22][24] = 8;
        pixel_data[22][25] = 9;
        pixel_data[22][26] = 9;
        pixel_data[22][27] = 9;
        pixel_data[22][28] = 9;
        pixel_data[22][29] = 9;
        pixel_data[22][30] = 9;
        pixel_data[22][31] = 9;
        pixel_data[22][32] = 9;
        pixel_data[22][33] = 9;
        pixel_data[22][34] = 10;
        pixel_data[22][35] = 10;
        pixel_data[22][36] = 6;
        pixel_data[22][37] = 6;
        pixel_data[22][38] = 6;
        pixel_data[22][39] = 6;
        pixel_data[22][40] = 11;
        pixel_data[22][41] = 1;
        pixel_data[22][42] = 11;
        pixel_data[22][43] = 11;
        pixel_data[22][44] = 11;
        pixel_data[22][45] = 11;
        pixel_data[22][46] = 11;
        pixel_data[22][47] = 11;
        pixel_data[22][48] = 11;
        pixel_data[22][49] = 11; // y=22
        pixel_data[23][0] = 1;
        pixel_data[23][1] = 1;
        pixel_data[23][2] = 1;
        pixel_data[23][3] = 1;
        pixel_data[23][4] = 1;
        pixel_data[23][5] = 12;
        pixel_data[23][6] = 6;
        pixel_data[23][7] = 7;
        pixel_data[23][8] = 7;
        pixel_data[23][9] = 10;
        pixel_data[23][10] = 8;
        pixel_data[23][11] = 9;
        pixel_data[23][12] = 9;
        pixel_data[23][13] = 9;
        pixel_data[23][14] = 9;
        pixel_data[23][15] = 9;
        pixel_data[23][16] = 9;
        pixel_data[23][17] = 10;
        pixel_data[23][18] = 10;
        pixel_data[23][19] = 6;
        pixel_data[23][20] = 6;
        pixel_data[23][21] = 6;
        pixel_data[23][22] = 6;
        pixel_data[23][23] = 6;
        pixel_data[23][24] = 8;
        pixel_data[23][25] = 9;
        pixel_data[23][26] = 9;
        pixel_data[23][27] = 9;
        pixel_data[23][28] = 9;
        pixel_data[23][29] = 9;
        pixel_data[23][30] = 9;
        pixel_data[23][31] = 9;
        pixel_data[23][32] = 9;
        pixel_data[23][33] = 9;
        pixel_data[23][34] = 8;
        pixel_data[23][35] = 10;
        pixel_data[23][36] = 6;
        pixel_data[23][37] = 6;
        pixel_data[23][38] = 6;
        pixel_data[23][39] = 6;
        pixel_data[23][40] = 7;
        pixel_data[23][41] = 11;
        pixel_data[23][42] = 11;
        pixel_data[23][43] = 11;
        pixel_data[23][44] = 11;
        pixel_data[23][45] = 11;
        pixel_data[23][46] = 11;
        pixel_data[23][47] = 11;
        pixel_data[23][48] = 11;
        pixel_data[23][49] = 11; // y=23
        pixel_data[24][0] = 1;
        pixel_data[24][1] = 1;
        pixel_data[24][2] = 1;
        pixel_data[24][3] = 1;
        pixel_data[24][4] = 1;
        pixel_data[24][5] = 7;
        pixel_data[24][6] = 6;
        pixel_data[24][7] = 6;
        pixel_data[24][8] = 7;
        pixel_data[24][9] = 10;
        pixel_data[24][10] = 8;
        pixel_data[24][11] = 9;
        pixel_data[24][12] = 9;
        pixel_data[24][13] = 9;
        pixel_data[24][14] = 9;
        pixel_data[24][15] = 9;
        pixel_data[24][16] = 8;
        pixel_data[24][17] = 10;
        pixel_data[24][18] = 7;
        pixel_data[24][19] = 6;
        pixel_data[24][20] = 6;
        pixel_data[24][21] = 6;
        pixel_data[24][22] = 6;
        pixel_data[24][23] = 6;
        pixel_data[24][24] = 8;
        pixel_data[24][25] = 9;
        pixel_data[24][26] = 9;
        pixel_data[24][27] = 9;
        pixel_data[24][28] = 9;
        pixel_data[24][29] = 9;
        pixel_data[24][30] = 9;
        pixel_data[24][31] = 9;
        pixel_data[24][32] = 9;
        pixel_data[24][33] = 9;
        pixel_data[24][34] = 8;
        pixel_data[24][35] = 10;
        pixel_data[24][36] = 6;
        pixel_data[24][37] = 6;
        pixel_data[24][38] = 6;
        pixel_data[24][39] = 6;
        pixel_data[24][40] = 6;
        pixel_data[24][41] = 7;
        pixel_data[24][42] = 1;
        pixel_data[24][43] = 11;
        pixel_data[24][44] = 11;
        pixel_data[24][45] = 11;
        pixel_data[24][46] = 11;
        pixel_data[24][47] = 11;
        pixel_data[24][48] = 11;
        pixel_data[24][49] = 11; // y=24
        pixel_data[25][0] = 1;
        pixel_data[25][1] = 1;
        pixel_data[25][2] = 1;
        pixel_data[25][3] = 1;
        pixel_data[25][4] = 1;
        pixel_data[25][5] = 7;
        pixel_data[25][6] = 6;
        pixel_data[25][7] = 6;
        pixel_data[25][8] = 7;
        pixel_data[25][9] = 10;
        pixel_data[25][10] = 8;
        pixel_data[25][11] = 9;
        pixel_data[25][12] = 9;
        pixel_data[25][13] = 9;
        pixel_data[25][14] = 9;
        pixel_data[25][15] = 8;
        pixel_data[25][16] = 10;
        pixel_data[25][17] = 10;
        pixel_data[25][18] = 6;
        pixel_data[25][19] = 6;
        pixel_data[25][20] = 6;
        pixel_data[25][21] = 6;
        pixel_data[25][22] = 6;
        pixel_data[25][23] = 10;
        pixel_data[25][24] = 8;
        pixel_data[25][25] = 9;
        pixel_data[25][26] = 9;
        pixel_data[25][27] = 9;
        pixel_data[25][28] = 9;
        pixel_data[25][29] = 9;
        pixel_data[25][30] = 9;
        pixel_data[25][31] = 9;
        pixel_data[25][32] = 9;
        pixel_data[25][33] = 9;
        pixel_data[25][34] = 8;
        pixel_data[25][35] = 10;
        pixel_data[25][36] = 7;
        pixel_data[25][37] = 6;
        pixel_data[25][38] = 6;
        pixel_data[25][39] = 6;
        pixel_data[25][40] = 6;
        pixel_data[25][41] = 6;
        pixel_data[25][42] = 11;
        pixel_data[25][43] = 1;
        pixel_data[25][44] = 11;
        pixel_data[25][45] = 11;
        pixel_data[25][46] = 11;
        pixel_data[25][47] = 11;
        pixel_data[25][48] = 11;
        pixel_data[25][49] = 11; // y=25
        pixel_data[26][0] = 11;
        pixel_data[26][1] = 1;
        pixel_data[26][2] = 1;
        pixel_data[26][3] = 1;
        pixel_data[26][4] = 11;
        pixel_data[26][5] = 7;
        pixel_data[26][6] = 7;
        pixel_data[26][7] = 6;
        pixel_data[26][8] = 6;
        pixel_data[26][9] = 10;
        pixel_data[26][10] = 10;
        pixel_data[26][11] = 9;
        pixel_data[26][12] = 9;
        pixel_data[26][13] = 9;
        pixel_data[26][14] = 9;
        pixel_data[26][15] = 10;
        pixel_data[26][16] = 10;
        pixel_data[26][17] = 6;
        pixel_data[26][18] = 6;
        pixel_data[26][19] = 6;
        pixel_data[26][20] = 6;
        pixel_data[26][21] = 6;
        pixel_data[26][22] = 7;
        pixel_data[26][23] = 10;
        pixel_data[26][24] = 10;
        pixel_data[26][25] = 9;
        pixel_data[26][26] = 9;
        pixel_data[26][27] = 9;
        pixel_data[26][28] = 9;
        pixel_data[26][29] = 9;
        pixel_data[26][30] = 9;
        pixel_data[26][31] = 9;
        pixel_data[26][32] = 9;
        pixel_data[26][33] = 9;
        pixel_data[26][34] = 10;
        pixel_data[26][35] = 10;
        pixel_data[26][36] = 6;
        pixel_data[26][37] = 6;
        pixel_data[26][38] = 6;
        pixel_data[26][39] = 6;
        pixel_data[26][40] = 6;
        pixel_data[26][41] = 6;
        pixel_data[26][42] = 7;
        pixel_data[26][43] = 11;
        pixel_data[26][44] = 1;
        pixel_data[26][45] = 11;
        pixel_data[26][46] = 11;
        pixel_data[26][47] = 11;
        pixel_data[26][48] = 11;
        pixel_data[26][49] = 11; // y=26
        pixel_data[27][0] = 11;
        pixel_data[27][1] = 1;
        pixel_data[27][2] = 1;
        pixel_data[27][3] = 1;
        pixel_data[27][4] = 7;
        pixel_data[27][5] = 7;
        pixel_data[27][6] = 7;
        pixel_data[27][7] = 6;
        pixel_data[27][8] = 6;
        pixel_data[27][9] = 10;
        pixel_data[27][10] = 10;
        pixel_data[27][11] = 10;
        pixel_data[27][12] = 9;
        pixel_data[27][13] = 8;
        pixel_data[27][14] = 10;
        pixel_data[27][15] = 10;
        pixel_data[27][16] = 7;
        pixel_data[27][17] = 6;
        pixel_data[27][18] = 6;
        pixel_data[27][19] = 6;
        pixel_data[27][20] = 6;
        pixel_data[27][21] = 6;
        pixel_data[27][22] = 6;
        pixel_data[27][23] = 10;
        pixel_data[27][24] = 10;
        pixel_data[27][25] = 8;
        pixel_data[27][26] = 9;
        pixel_data[27][27] = 9;
        pixel_data[27][28] = 9;
        pixel_data[27][29] = 9;
        pixel_data[27][30] = 9;
        pixel_data[27][31] = 9;
        pixel_data[27][32] = 9;
        pixel_data[27][33] = 8;
        pixel_data[27][34] = 10;
        pixel_data[27][35] = 10;
        pixel_data[27][36] = 6;
        pixel_data[27][37] = 6;
        pixel_data[27][38] = 6;
        pixel_data[27][39] = 6;
        pixel_data[27][40] = 6;
        pixel_data[27][41] = 6;
        pixel_data[27][42] = 6;
        pixel_data[27][43] = 7;
        pixel_data[27][44] = 1;
        pixel_data[27][45] = 11;
        pixel_data[27][46] = 11;
        pixel_data[27][47] = 11;
        pixel_data[27][48] = 11;
        pixel_data[27][49] = 11; // y=27
        pixel_data[28][0] = 11;
        pixel_data[28][1] = 1;
        pixel_data[28][2] = 1;
        pixel_data[28][3] = 12;
        pixel_data[28][4] = 7;
        pixel_data[28][5] = 7;
        pixel_data[28][6] = 7;
        pixel_data[28][7] = 6;
        pixel_data[28][8] = 6;
        pixel_data[28][9] = 10;
        pixel_data[28][10] = 10;
        pixel_data[28][11] = 10;
        pixel_data[28][12] = 10;
        pixel_data[28][13] = 10;
        pixel_data[28][14] = 10;
        pixel_data[28][15] = 10;
        pixel_data[28][16] = 6;
        pixel_data[28][17] = 6;
        pixel_data[28][18] = 6;
        pixel_data[28][19] = 6;
        pixel_data[28][20] = 6;
        pixel_data[28][21] = 6;
        pixel_data[28][22] = 6;
        pixel_data[28][23] = 10;
        pixel_data[28][24] = 10;
        pixel_data[28][25] = 10;
        pixel_data[28][26] = 9;
        pixel_data[28][27] = 9;
        pixel_data[28][28] = 9;
        pixel_data[28][29] = 9;
        pixel_data[28][30] = 9;
        pixel_data[28][31] = 8;
        pixel_data[28][32] = 10;
        pixel_data[28][33] = 10;
        pixel_data[28][34] = 10;
        pixel_data[28][35] = 7;
        pixel_data[28][36] = 6;
        pixel_data[28][37] = 6;
        pixel_data[28][38] = 6;
        pixel_data[28][39] = 6;
        pixel_data[28][40] = 6;
        pixel_data[28][41] = 6;
        pixel_data[28][42] = 6;
        pixel_data[28][43] = 6;
        pixel_data[28][44] = 11;
        pixel_data[28][45] = 1;
        pixel_data[28][46] = 11;
        pixel_data[28][47] = 11;
        pixel_data[28][48] = 11;
        pixel_data[28][49] = 0; // y=28
        pixel_data[29][0] = 11;
        pixel_data[29][1] = 1;
        pixel_data[29][2] = 1;
        pixel_data[29][3] = 7;
        pixel_data[29][4] = 7;
        pixel_data[29][5] = 7;
        pixel_data[29][6] = 7;
        pixel_data[29][7] = 6;
        pixel_data[29][8] = 6;
        pixel_data[29][9] = 6;
        pixel_data[29][10] = 7;
        pixel_data[29][11] = 10;
        pixel_data[29][12] = 10;
        pixel_data[29][13] = 10;
        pixel_data[29][14] = 10;
        pixel_data[29][15] = 6;
        pixel_data[29][16] = 6;
        pixel_data[29][17] = 6;
        pixel_data[29][18] = 6;
        pixel_data[29][19] = 6;
        pixel_data[29][20] = 6;
        pixel_data[29][21] = 6;
        pixel_data[29][22] = 6;
        pixel_data[29][23] = 6;
        pixel_data[29][24] = 10;
        pixel_data[29][25] = 10;
        pixel_data[29][26] = 10;
        pixel_data[29][27] = 8;
        pixel_data[29][28] = 9;
        pixel_data[29][29] = 9;
        pixel_data[29][30] = 8;
        pixel_data[29][31] = 10;
        pixel_data[29][32] = 10;
        pixel_data[29][33] = 10;
        pixel_data[29][34] = 10;
        pixel_data[29][35] = 6;
        pixel_data[29][36] = 6;
        pixel_data[29][37] = 6;
        pixel_data[29][38] = 6;
        pixel_data[29][39] = 6;
        pixel_data[29][40] = 6;
        pixel_data[29][41] = 6;
        pixel_data[29][42] = 6;
        pixel_data[29][43] = 6;
        pixel_data[29][44] = 7;
        pixel_data[29][45] = 1;
        pixel_data[29][46] = 11;
        pixel_data[29][47] = 11;
        pixel_data[29][48] = 11;
        pixel_data[29][49] = 0; // y=29
        pixel_data[30][0] = 7;
        pixel_data[30][1] = 1;
        pixel_data[30][2] = 1;
        pixel_data[30][3] = 7;
        pixel_data[30][4] = 7;
        pixel_data[30][5] = 7;
        pixel_data[30][6] = 7;
        pixel_data[30][7] = 6;
        pixel_data[30][8] = 6;
        pixel_data[30][9] = 6;
        pixel_data[30][10] = 6;
        pixel_data[30][11] = 6;
        pixel_data[30][12] = 7;
        pixel_data[30][13] = 6;
        pixel_data[30][14] = 6;
        pixel_data[30][15] = 6;
        pixel_data[30][16] = 6;
        pixel_data[30][17] = 6;
        pixel_data[30][18] = 6;
        pixel_data[30][19] = 6;
        pixel_data[30][20] = 6;
        pixel_data[30][21] = 6;
        pixel_data[30][22] = 6;
        pixel_data[30][23] = 6;
        pixel_data[30][24] = 7;
        pixel_data[30][25] = 10;
        pixel_data[30][26] = 10;
        pixel_data[30][27] = 10;
        pixel_data[30][28] = 10;
        pixel_data[30][29] = 10;
        pixel_data[30][30] = 10;
        pixel_data[30][31] = 10;
        pixel_data[30][32] = 10;
        pixel_data[30][33] = 10;
        pixel_data[30][34] = 6;
        pixel_data[30][35] = 6;
        pixel_data[30][36] = 6;
        pixel_data[30][37] = 6;
        pixel_data[30][38] = 6;
        pixel_data[30][39] = 6;
        pixel_data[30][40] = 6;
        pixel_data[30][41] = 6;
        pixel_data[30][42] = 6;
        pixel_data[30][43] = 6;
        pixel_data[30][44] = 6;
        pixel_data[30][45] = 11;
        pixel_data[30][46] = 1;
        pixel_data[30][47] = 11;
        pixel_data[30][48] = 11;
        pixel_data[30][49] = 0; // y=30
        pixel_data[31][0] = 0;
        pixel_data[31][1] = 1;
        pixel_data[31][2] = 11;
        pixel_data[31][3] = 7;
        pixel_data[31][4] = 7;
        pixel_data[31][5] = 7;
        pixel_data[31][6] = 6;
        pixel_data[31][7] = 6;
        pixel_data[31][8] = 6;
        pixel_data[31][9] = 6;
        pixel_data[31][10] = 6;
        pixel_data[31][11] = 6;
        pixel_data[31][12] = 6;
        pixel_data[31][13] = 6;
        pixel_data[31][14] = 7;
        pixel_data[31][15] = 7;
        pixel_data[31][16] = 7;
        pixel_data[31][17] = 7;
        pixel_data[31][18] = 7;
        pixel_data[31][19] = 6;
        pixel_data[31][20] = 6;
        pixel_data[31][21] = 6;
        pixel_data[31][22] = 6;
        pixel_data[31][23] = 6;
        pixel_data[31][24] = 6;
        pixel_data[31][25] = 6;
        pixel_data[31][26] = 7;
        pixel_data[31][27] = 10;
        pixel_data[31][28] = 10;
        pixel_data[31][29] = 10;
        pixel_data[31][30] = 10;
        pixel_data[31][31] = 10;
        pixel_data[31][32] = 7;
        pixel_data[31][33] = 6;
        pixel_data[31][34] = 6;
        pixel_data[31][35] = 6;
        pixel_data[31][36] = 6;
        pixel_data[31][37] = 6;
        pixel_data[31][38] = 6;
        pixel_data[31][39] = 6;
        pixel_data[31][40] = 6;
        pixel_data[31][41] = 6;
        pixel_data[31][42] = 6;
        pixel_data[31][43] = 6;
        pixel_data[31][44] = 6;
        pixel_data[31][45] = 7;
        pixel_data[31][46] = 11;
        pixel_data[31][47] = 11;
        pixel_data[31][48] = 0;
        pixel_data[31][49] = 1; // y=31
        pixel_data[32][0] = 0;
        pixel_data[32][1] = 1;
        pixel_data[32][2] = 7;
        pixel_data[32][3] = 6;
        pixel_data[32][4] = 6;
        pixel_data[32][5] = 6;
        pixel_data[32][6] = 6;
        pixel_data[32][7] = 6;
        pixel_data[32][8] = 6;
        pixel_data[32][9] = 6;
        pixel_data[32][10] = 6;
        pixel_data[32][11] = 7;
        pixel_data[32][12] = 10;
        pixel_data[32][13] = 10;
        pixel_data[32][14] = 10;
        pixel_data[32][15] = 10;
        pixel_data[32][16] = 10;
        pixel_data[32][17] = 10;
        pixel_data[32][18] = 10;
        pixel_data[32][19] = 10;
        pixel_data[32][20] = 10;
        pixel_data[32][21] = 10;
        pixel_data[32][22] = 7;
        pixel_data[32][23] = 6;
        pixel_data[32][24] = 6;
        pixel_data[32][25] = 6;
        pixel_data[32][26] = 6;
        pixel_data[32][27] = 6;
        pixel_data[32][28] = 6;
        pixel_data[32][29] = 6;
        pixel_data[32][30] = 6;
        pixel_data[32][31] = 6;
        pixel_data[32][32] = 6;
        pixel_data[32][33] = 6;
        pixel_data[32][34] = 6;
        pixel_data[32][35] = 6;
        pixel_data[32][36] = 6;
        pixel_data[32][37] = 6;
        pixel_data[32][38] = 6;
        pixel_data[32][39] = 6;
        pixel_data[32][40] = 6;
        pixel_data[32][41] = 6;
        pixel_data[32][42] = 6;
        pixel_data[32][43] = 6;
        pixel_data[32][44] = 6;
        pixel_data[32][45] = 6;
        pixel_data[32][46] = 11;
        pixel_data[32][47] = 1;
        pixel_data[32][48] = 0;
        pixel_data[32][49] = 5; // y=32
        pixel_data[33][0] = 0;
        pixel_data[33][1] = 6;
        pixel_data[33][2] = 6;
        pixel_data[33][3] = 6;
        pixel_data[33][4] = 6;
        pixel_data[33][5] = 6;
        pixel_data[33][6] = 6;
        pixel_data[33][7] = 6;
        pixel_data[33][8] = 6;
        pixel_data[33][9] = 7;
        pixel_data[33][10] = 10;
        pixel_data[33][11] = 10;
        pixel_data[33][12] = 10;
        pixel_data[33][13] = 10;
        pixel_data[33][14] = 10;
        pixel_data[33][15] = 10;
        pixel_data[33][16] = 7;
        pixel_data[33][17] = 7;
        pixel_data[33][18] = 10;
        pixel_data[33][19] = 10;
        pixel_data[33][20] = 10;
        pixel_data[33][21] = 10;
        pixel_data[33][22] = 10;
        pixel_data[33][23] = 10;
        pixel_data[33][24] = 7;
        pixel_data[33][25] = 6;
        pixel_data[33][26] = 6;
        pixel_data[33][27] = 6;
        pixel_data[33][28] = 6;
        pixel_data[33][29] = 6;
        pixel_data[33][30] = 6;
        pixel_data[33][31] = 6;
        pixel_data[33][32] = 6;
        pixel_data[33][33] = 6;
        pixel_data[33][34] = 6;
        pixel_data[33][35] = 6;
        pixel_data[33][36] = 6;
        pixel_data[33][37] = 6;
        pixel_data[33][38] = 6;
        pixel_data[33][39] = 6;
        pixel_data[33][40] = 6;
        pixel_data[33][41] = 6;
        pixel_data[33][42] = 6;
        pixel_data[33][43] = 6;
        pixel_data[33][44] = 6;
        pixel_data[33][45] = 6;
        pixel_data[33][46] = 7;
        pixel_data[33][47] = 1;
        pixel_data[33][48] = 0;
        pixel_data[33][49] = 1; // y=33
        pixel_data[34][0] = 0;
        pixel_data[34][1] = 14;
        pixel_data[34][2] = 4;
        pixel_data[34][3] = 7;
        pixel_data[34][4] = 6;
        pixel_data[34][5] = 6;
        pixel_data[34][6] = 6;
        pixel_data[34][7] = 6;
        pixel_data[34][8] = 10;
        pixel_data[34][9] = 10;
        pixel_data[34][10] = 10;
        pixel_data[34][11] = 10;
        pixel_data[34][12] = 6;
        pixel_data[34][13] = 6;
        pixel_data[34][14] = 6;
        pixel_data[34][15] = 6;
        pixel_data[34][16] = 6;
        pixel_data[34][17] = 6;
        pixel_data[34][18] = 6;
        pixel_data[34][19] = 6;
        pixel_data[34][20] = 6;
        pixel_data[34][21] = 7;
        pixel_data[34][22] = 10;
        pixel_data[34][23] = 10;
        pixel_data[34][24] = 10;
        pixel_data[34][25] = 10;
        pixel_data[34][26] = 7;
        pixel_data[34][27] = 6;
        pixel_data[34][28] = 6;
        pixel_data[34][29] = 6;
        pixel_data[34][30] = 6;
        pixel_data[34][31] = 6;
        pixel_data[34][32] = 6;
        pixel_data[34][33] = 6;
        pixel_data[34][34] = 6;
        pixel_data[34][35] = 6;
        pixel_data[34][36] = 6;
        pixel_data[34][37] = 6;
        pixel_data[34][38] = 6;
        pixel_data[34][39] = 6;
        pixel_data[34][40] = 6;
        pixel_data[34][41] = 6;
        pixel_data[34][42] = 6;
        pixel_data[34][43] = 6;
        pixel_data[34][44] = 6;
        pixel_data[34][45] = 6;
        pixel_data[34][46] = 15;
        pixel_data[34][47] = 14;
        pixel_data[34][48] = 0;
        pixel_data[34][49] = 12; // y=34
        pixel_data[35][0] = 0;
        pixel_data[35][1] = 13;
        pixel_data[35][2] = 15;
        pixel_data[35][3] = 6;
        pixel_data[35][4] = 6;
        pixel_data[35][5] = 6;
        pixel_data[35][6] = 6;
        pixel_data[35][7] = 10;
        pixel_data[35][8] = 10;
        pixel_data[35][9] = 10;
        pixel_data[35][10] = 6;
        pixel_data[35][11] = 6;
        pixel_data[35][12] = 6;
        pixel_data[35][13] = 6;
        pixel_data[35][14] = 6;
        pixel_data[35][15] = 6;
        pixel_data[35][16] = 6;
        pixel_data[35][17] = 6;
        pixel_data[35][18] = 6;
        pixel_data[35][19] = 6;
        pixel_data[35][20] = 6;
        pixel_data[35][21] = 6;
        pixel_data[35][22] = 6;
        pixel_data[35][23] = 6;
        pixel_data[35][24] = 10;
        pixel_data[35][25] = 10;
        pixel_data[35][26] = 10;
        pixel_data[35][27] = 10;
        pixel_data[35][28] = 6;
        pixel_data[35][29] = 6;
        pixel_data[35][30] = 6;
        pixel_data[35][31] = 6;
        pixel_data[35][32] = 6;
        pixel_data[35][33] = 6;
        pixel_data[35][34] = 6;
        pixel_data[35][35] = 6;
        pixel_data[35][36] = 6;
        pixel_data[35][37] = 6;
        pixel_data[35][38] = 6;
        pixel_data[35][39] = 6;
        pixel_data[35][40] = 6;
        pixel_data[35][41] = 6;
        pixel_data[35][42] = 6;
        pixel_data[35][43] = 6;
        pixel_data[35][44] = 7;
        pixel_data[35][45] = 6;
        pixel_data[35][46] = 13;
        pixel_data[35][47] = 13;
        pixel_data[35][48] = 0;
        pixel_data[35][49] = 14; // y=35
        pixel_data[36][0] = 0;
        pixel_data[36][1] = 13;
        pixel_data[36][2] = 12;
        pixel_data[36][3] = 4;
        pixel_data[36][4] = 7;
        pixel_data[36][5] = 6;
        pixel_data[36][6] = 10;
        pixel_data[36][7] = 10;
        pixel_data[36][8] = 10;
        pixel_data[36][9] = 6;
        pixel_data[36][10] = 6;
        pixel_data[36][11] = 6;
        pixel_data[36][12] = 6;
        pixel_data[36][13] = 6;
        pixel_data[36][14] = 6;
        pixel_data[36][15] = 6;
        pixel_data[36][16] = 6;
        pixel_data[36][17] = 6;
        pixel_data[36][18] = 6;
        pixel_data[36][19] = 6;
        pixel_data[36][20] = 6;
        pixel_data[36][21] = 6;
        pixel_data[36][22] = 6;
        pixel_data[36][23] = 6;
        pixel_data[36][24] = 6;
        pixel_data[36][25] = 7;
        pixel_data[36][26] = 10;
        pixel_data[36][27] = 10;
        pixel_data[36][28] = 10;
        pixel_data[36][29] = 6;
        pixel_data[36][30] = 6;
        pixel_data[36][31] = 6;
        pixel_data[36][32] = 6;
        pixel_data[36][33] = 6;
        pixel_data[36][34] = 6;
        pixel_data[36][35] = 6;
        pixel_data[36][36] = 6;
        pixel_data[36][37] = 6;
        pixel_data[36][38] = 6;
        pixel_data[36][39] = 6;
        pixel_data[36][40] = 6;
        pixel_data[36][41] = 6;
        pixel_data[36][42] = 6;
        pixel_data[36][43] = 6;
        pixel_data[36][44] = 6;
        pixel_data[36][45] = 15;
        pixel_data[36][46] = 13;
        pixel_data[36][47] = 3;
        pixel_data[36][48] = 0;
        pixel_data[36][49] = 15; // y=36
        pixel_data[37][0] = 0;
        pixel_data[37][1] = 13;
        pixel_data[37][2] = 13;
        pixel_data[37][3] = 3;
        pixel_data[37][4] = 6;
        pixel_data[37][5] = 7;
        pixel_data[37][6] = 10;
        pixel_data[37][7] = 10;
        pixel_data[37][8] = 6;
        pixel_data[37][9] = 6;
        pixel_data[37][10] = 6;
        pixel_data[37][11] = 6;
        pixel_data[37][12] = 6;
        pixel_data[37][13] = 6;
        pixel_data[37][14] = 6;
        pixel_data[37][15] = 6;
        pixel_data[37][16] = 6;
        pixel_data[37][17] = 6;
        pixel_data[37][18] = 6;
        pixel_data[37][19] = 6;
        pixel_data[37][20] = 6;
        pixel_data[37][21] = 6;
        pixel_data[37][22] = 6;
        pixel_data[37][23] = 6;
        pixel_data[37][24] = 6;
        pixel_data[37][25] = 6;
        pixel_data[37][26] = 6;
        pixel_data[37][27] = 10;
        pixel_data[37][28] = 10;
        pixel_data[37][29] = 10;
        pixel_data[37][30] = 6;
        pixel_data[37][31] = 6;
        pixel_data[37][32] = 6;
        pixel_data[37][33] = 6;
        pixel_data[37][34] = 6;
        pixel_data[37][35] = 6;
        pixel_data[37][36] = 6;
        pixel_data[37][37] = 6;
        pixel_data[37][38] = 6;
        pixel_data[37][39] = 6;
        pixel_data[37][40] = 6;
        pixel_data[37][41] = 6;
        pixel_data[37][42] = 6;
        pixel_data[37][43] = 7;
        pixel_data[37][44] = 4;
        pixel_data[37][45] = 13;
        pixel_data[37][46] = 13;
        pixel_data[37][47] = 13;
        pixel_data[37][48] = 0;
        pixel_data[37][49] = 15; // y=37
        pixel_data[38][0] = 0;
        pixel_data[38][1] = 13;
        pixel_data[38][2] = 13;
        pixel_data[38][3] = 13;
        pixel_data[38][4] = 15;
        pixel_data[38][5] = 7;
        pixel_data[38][6] = 10;
        pixel_data[38][7] = 6;
        pixel_data[38][8] = 6;
        pixel_data[38][9] = 6;
        pixel_data[38][10] = 6;
        pixel_data[38][11] = 6;
        pixel_data[38][12] = 6;
        pixel_data[38][13] = 6;
        pixel_data[38][14] = 6;
        pixel_data[38][15] = 6;
        pixel_data[38][16] = 6;
        pixel_data[38][17] = 6;
        pixel_data[38][18] = 6;
        pixel_data[38][19] = 6;
        pixel_data[38][20] = 6;
        pixel_data[38][21] = 6;
        pixel_data[38][22] = 6;
        pixel_data[38][23] = 6;
        pixel_data[38][24] = 6;
        pixel_data[38][25] = 6;
        pixel_data[38][26] = 6;
        pixel_data[38][27] = 6;
        pixel_data[38][28] = 10;
        pixel_data[38][29] = 10;
        pixel_data[38][30] = 10;
        pixel_data[38][31] = 6;
        pixel_data[38][32] = 6;
        pixel_data[38][33] = 6;
        pixel_data[38][34] = 6;
        pixel_data[38][35] = 6;
        pixel_data[38][36] = 6;
        pixel_data[38][37] = 6;
        pixel_data[38][38] = 6;
        pixel_data[38][39] = 6;
        pixel_data[38][40] = 6;
        pixel_data[38][41] = 6;
        pixel_data[38][42] = 7;
        pixel_data[38][43] = 4;
        pixel_data[38][44] = 13;
        pixel_data[38][45] = 13;
        pixel_data[38][46] = 13;
        pixel_data[38][47] = 13;
        pixel_data[38][48] = 0;
        pixel_data[38][49] = 15; // y=38
        pixel_data[39][0] = 0;
        pixel_data[39][1] = 13;
        pixel_data[39][2] = 13;
        pixel_data[39][3] = 13;
        pixel_data[39][4] = 13;
        pixel_data[39][5] = 4;
        pixel_data[39][6] = 7;
        pixel_data[39][7] = 6;
        pixel_data[39][8] = 6;
        pixel_data[39][9] = 6;
        pixel_data[39][10] = 6;
        pixel_data[39][11] = 6;
        pixel_data[39][12] = 6;
        pixel_data[39][13] = 6;
        pixel_data[39][14] = 6;
        pixel_data[39][15] = 6;
        pixel_data[39][16] = 6;
        pixel_data[39][17] = 6;
        pixel_data[39][18] = 6;
        pixel_data[39][19] = 6;
        pixel_data[39][20] = 6;
        pixel_data[39][21] = 6;
        pixel_data[39][22] = 6;
        pixel_data[39][23] = 6;
        pixel_data[39][24] = 6;
        pixel_data[39][25] = 6;
        pixel_data[39][26] = 6;
        pixel_data[39][27] = 6;
        pixel_data[39][28] = 6;
        pixel_data[39][29] = 10;
        pixel_data[39][30] = 10;
        pixel_data[39][31] = 7;
        pixel_data[39][32] = 6;
        pixel_data[39][33] = 6;
        pixel_data[39][34] = 6;
        pixel_data[39][35] = 6;
        pixel_data[39][36] = 6;
        pixel_data[39][37] = 6;
        pixel_data[39][38] = 6;
        pixel_data[39][39] = 6;
        pixel_data[39][40] = 6;
        pixel_data[39][41] = 7;
        pixel_data[39][42] = 6;
        pixel_data[39][43] = 13;
        pixel_data[39][44] = 13;
        pixel_data[39][45] = 13;
        pixel_data[39][46] = 13;
        pixel_data[39][47] = 13;
        pixel_data[39][48] = 0;
        pixel_data[39][49] = 15; // y=39
        pixel_data[40][0] = 0;
        pixel_data[40][1] = 13;
        pixel_data[40][2] = 13;
        pixel_data[40][3] = 13;
        pixel_data[40][4] = 13;
        pixel_data[40][5] = 13;
        pixel_data[40][6] = 4;
        pixel_data[40][7] = 7;
        pixel_data[40][8] = 6;
        pixel_data[40][9] = 6;
        pixel_data[40][10] = 6;
        pixel_data[40][11] = 6;
        pixel_data[40][12] = 6;
        pixel_data[40][13] = 6;
        pixel_data[40][14] = 6;
        pixel_data[40][15] = 6;
        pixel_data[40][16] = 6;
        pixel_data[40][17] = 6;
        pixel_data[40][18] = 6;
        pixel_data[40][19] = 6;
        pixel_data[40][20] = 6;
        pixel_data[40][21] = 6;
        pixel_data[40][22] = 6;
        pixel_data[40][23] = 6;
        pixel_data[40][24] = 6;
        pixel_data[40][25] = 6;
        pixel_data[40][26] = 6;
        pixel_data[40][27] = 6;
        pixel_data[40][28] = 6;
        pixel_data[40][29] = 6;
        pixel_data[40][30] = 10;
        pixel_data[40][31] = 10;
        pixel_data[40][32] = 6;
        pixel_data[40][33] = 6;
        pixel_data[40][34] = 6;
        pixel_data[40][35] = 6;
        pixel_data[40][36] = 6;
        pixel_data[40][37] = 6;
        pixel_data[40][38] = 6;
        pixel_data[40][39] = 6;
        pixel_data[40][40] = 7;
        pixel_data[40][41] = 6;
        pixel_data[40][42] = 3;
        pixel_data[40][43] = 13;
        pixel_data[40][44] = 13;
        pixel_data[40][45] = 13;
        pixel_data[40][46] = 13;
        pixel_data[40][47] = 13;
        pixel_data[40][48] = 0;
        pixel_data[40][49] = 4; // y=40
        pixel_data[41][0] = 0;
        pixel_data[41][1] = 13;
        pixel_data[41][2] = 13;
        pixel_data[41][3] = 13;
        pixel_data[41][4] = 13;
        pixel_data[41][5] = 13;
        pixel_data[41][6] = 13;
        pixel_data[41][7] = 4;
        pixel_data[41][8] = 7;
        pixel_data[41][9] = 6;
        pixel_data[41][10] = 6;
        pixel_data[41][11] = 6;
        pixel_data[41][12] = 6;
        pixel_data[41][13] = 6;
        pixel_data[41][14] = 6;
        pixel_data[41][15] = 6;
        pixel_data[41][16] = 6;
        pixel_data[41][17] = 6;
        pixel_data[41][18] = 6;
        pixel_data[41][19] = 6;
        pixel_data[41][20] = 6;
        pixel_data[41][21] = 6;
        pixel_data[41][22] = 6;
        pixel_data[41][23] = 6;
        pixel_data[41][24] = 6;
        pixel_data[41][25] = 6;
        pixel_data[41][26] = 6;
        pixel_data[41][27] = 6;
        pixel_data[41][28] = 6;
        pixel_data[41][29] = 6;
        pixel_data[41][30] = 7;
        pixel_data[41][31] = 10;
        pixel_data[41][32] = 10;
        pixel_data[41][33] = 6;
        pixel_data[41][34] = 6;
        pixel_data[41][35] = 6;
        pixel_data[41][36] = 6;
        pixel_data[41][37] = 6;
        pixel_data[41][38] = 6;
        pixel_data[41][39] = 7;
        pixel_data[41][40] = 4;
        pixel_data[41][41] = 3;
        pixel_data[41][42] = 13;
        pixel_data[41][43] = 13;
        pixel_data[41][44] = 13;
        pixel_data[41][45] = 13;
        pixel_data[41][46] = 13;
        pixel_data[41][47] = 15;
        pixel_data[41][48] = 0;
        pixel_data[41][49] = 12; // y=41
        pixel_data[42][0] = 0;
        pixel_data[42][1] = 3;
        pixel_data[42][2] = 13;
        pixel_data[42][3] = 13;
        pixel_data[42][4] = 13;
        pixel_data[42][5] = 13;
        pixel_data[42][6] = 13;
        pixel_data[42][7] = 13;
        pixel_data[42][8] = 4;
        pixel_data[42][9] = 7;
        pixel_data[42][10] = 6;
        pixel_data[42][11] = 6;
        pixel_data[42][12] = 6;
        pixel_data[42][13] = 6;
        pixel_data[42][14] = 6;
        pixel_data[42][15] = 6;
        pixel_data[42][16] = 6;
        pixel_data[42][17] = 6;
        pixel_data[42][18] = 6;
        pixel_data[42][19] = 6;
        pixel_data[42][20] = 6;
        pixel_data[42][21] = 6;
        pixel_data[42][22] = 6;
        pixel_data[42][23] = 6;
        pixel_data[42][24] = 6;
        pixel_data[42][25] = 6;
        pixel_data[42][26] = 6;
        pixel_data[42][27] = 6;
        pixel_data[42][28] = 6;
        pixel_data[42][29] = 6;
        pixel_data[42][30] = 6;
        pixel_data[42][31] = 10;
        pixel_data[42][32] = 10;
        pixel_data[42][33] = 6;
        pixel_data[42][34] = 6;
        pixel_data[42][35] = 6;
        pixel_data[42][36] = 6;
        pixel_data[42][37] = 7;
        pixel_data[42][38] = 7;
        pixel_data[42][39] = 4;
        pixel_data[42][40] = 13;
        pixel_data[42][41] = 13;
        pixel_data[42][42] = 13;
        pixel_data[42][43] = 13;
        pixel_data[42][44] = 13;
        pixel_data[42][45] = 13;
        pixel_data[42][46] = 13;
        pixel_data[42][47] = 0;
        pixel_data[42][48] = 14;
        pixel_data[42][49] = 0; // y=42
        pixel_data[43][0] = 14;
        pixel_data[43][1] = 14;
        pixel_data[43][2] = 13;
        pixel_data[43][3] = 13;
        pixel_data[43][4] = 13;
        pixel_data[43][5] = 13;
        pixel_data[43][6] = 13;
        pixel_data[43][7] = 13;
        pixel_data[43][8] = 13;
        pixel_data[43][9] = 15;
        pixel_data[43][10] = 6;
        pixel_data[43][11] = 6;
        pixel_data[43][12] = 6;
        pixel_data[43][13] = 6;
        pixel_data[43][14] = 6;
        pixel_data[43][15] = 6;
        pixel_data[43][16] = 6;
        pixel_data[43][17] = 6;
        pixel_data[43][18] = 6;
        pixel_data[43][19] = 6;
        pixel_data[43][20] = 6;
        pixel_data[43][21] = 6;
        pixel_data[43][22] = 6;
        pixel_data[43][23] = 6;
        pixel_data[43][24] = 6;
        pixel_data[43][25] = 6;
        pixel_data[43][26] = 6;
        pixel_data[43][27] = 6;
        pixel_data[43][28] = 7;
        pixel_data[43][29] = 7;
        pixel_data[43][30] = 6;
        pixel_data[43][31] = 7;
        pixel_data[43][32] = 10;
        pixel_data[43][33] = 7;
        pixel_data[43][34] = 6;
        pixel_data[43][35] = 6;
        pixel_data[43][36] = 7;
        pixel_data[43][37] = 6;
        pixel_data[43][38] = 15;
        pixel_data[43][39] = 13;
        pixel_data[43][40] = 13;
        pixel_data[43][41] = 13;
        pixel_data[43][42] = 13;
        pixel_data[43][43] = 13;
        pixel_data[43][44] = 13;
        pixel_data[43][45] = 13;
        pixel_data[43][46] = 3;
        pixel_data[43][47] = 0;
        pixel_data[43][48] = 14;
        pixel_data[43][49] = 0; // y=43
        pixel_data[44][0] = 12;
        pixel_data[44][1] = 7;
        pixel_data[44][2] = 14;
        pixel_data[44][3] = 13;
        pixel_data[44][4] = 13;
        pixel_data[44][5] = 13;
        pixel_data[44][6] = 13;
        pixel_data[44][7] = 13;
        pixel_data[44][8] = 13;
        pixel_data[44][9] = 13;
        pixel_data[44][10] = 13;
        pixel_data[44][11] = 6;
        pixel_data[44][12] = 11;
        pixel_data[44][13] = 7;
        pixel_data[44][14] = 6;
        pixel_data[44][15] = 6;
        pixel_data[44][16] = 6;
        pixel_data[44][17] = 6;
        pixel_data[44][18] = 6;
        pixel_data[44][19] = 6;
        pixel_data[44][20] = 6;
        pixel_data[44][21] = 6;
        pixel_data[44][22] = 6;
        pixel_data[44][23] = 6;
        pixel_data[44][24] = 6;
        pixel_data[44][25] = 6;
        pixel_data[44][26] = 6;
        pixel_data[44][27] = 7;
        pixel_data[44][28] = 11;
        pixel_data[44][29] = 7;
        pixel_data[44][30] = 6;
        pixel_data[44][31] = 6;
        pixel_data[44][32] = 6;
        pixel_data[44][33] = 6;
        pixel_data[44][34] = 7;
        pixel_data[44][35] = 6;
        pixel_data[44][36] = 4;
        pixel_data[44][37] = 3;
        pixel_data[44][38] = 13;
        pixel_data[44][39] = 13;
        pixel_data[44][40] = 13;
        pixel_data[44][41] = 13;
        pixel_data[44][42] = 13;
        pixel_data[44][43] = 13;
        pixel_data[44][44] = 13;
        pixel_data[44][45] = 3;
        pixel_data[44][46] = 0;
        pixel_data[44][47] = 3;
        pixel_data[44][48] = 0;
        pixel_data[44][49] = 0; // y=44
        pixel_data[45][0] = 0;
        pixel_data[45][1] = 7;
        pixel_data[45][2] = 0;
        pixel_data[45][3] = 0;
        pixel_data[45][4] = 13;
        pixel_data[45][5] = 13;
        pixel_data[45][6] = 13;
        pixel_data[45][7] = 13;
        pixel_data[45][8] = 13;
        pixel_data[45][9] = 13;
        pixel_data[45][10] = 13;
        pixel_data[45][11] = 14;
        pixel_data[45][12] = 1;
        pixel_data[45][13] = 6;
        pixel_data[45][14] = 6;
        pixel_data[45][15] = 7;
        pixel_data[45][16] = 7;
        pixel_data[45][17] = 6;
        pixel_data[45][18] = 6;
        pixel_data[45][19] = 6;
        pixel_data[45][20] = 6;
        pixel_data[45][21] = 6;
        pixel_data[45][22] = 6;
        pixel_data[45][23] = 6;
        pixel_data[45][24] = 6;
        pixel_data[45][25] = 6;
        pixel_data[45][26] = 6;
        pixel_data[45][27] = 11;
        pixel_data[45][28] = 1;
        pixel_data[45][29] = 11;
        pixel_data[45][30] = 6;
        pixel_data[45][31] = 4;
        pixel_data[45][32] = 15;
        pixel_data[45][33] = 4;
        pixel_data[45][34] = 4;
        pixel_data[45][35] = 15;
        pixel_data[45][36] = 13;
        pixel_data[45][37] = 13;
        pixel_data[45][38] = 13;
        pixel_data[45][39] = 13;
        pixel_data[45][40] = 13;
        pixel_data[45][41] = 13;
        pixel_data[45][42] = 13;
        pixel_data[45][43] = 13;
        pixel_data[45][44] = 13;
        pixel_data[45][45] = 14;
        pixel_data[45][46] = 3;
        pixel_data[45][47] = 12;
        pixel_data[45][48] = 0;
        pixel_data[45][49] = 0; // y=45
        pixel_data[46][0] = 0;
        pixel_data[46][1] = 0;
        pixel_data[46][2] = 12;
        pixel_data[46][3] = 3;
        pixel_data[46][4] = 0;
        pixel_data[46][5] = 0;
        pixel_data[46][6] = 13;
        pixel_data[46][7] = 13;
        pixel_data[46][8] = 13;
        pixel_data[46][9] = 13;
        pixel_data[46][10] = 0;
        pixel_data[46][11] = 0;
        pixel_data[46][12] = 0;
        pixel_data[46][13] = 13;
        pixel_data[46][14] = 15;
        pixel_data[46][15] = 4;
        pixel_data[46][16] = 6;
        pixel_data[46][17] = 6;
        pixel_data[46][18] = 7;
        pixel_data[46][19] = 7;
        pixel_data[46][20] = 7;
        pixel_data[46][21] = 7;
        pixel_data[46][22] = 6;
        pixel_data[46][23] = 6;
        pixel_data[46][24] = 6;
        pixel_data[46][25] = 6;
        pixel_data[46][26] = 11;
        pixel_data[46][27] = 1;
        pixel_data[46][28] = 11;
        pixel_data[46][29] = 1;
        pixel_data[46][30] = 7;
        pixel_data[46][31] = 15;
        pixel_data[46][32] = 13;
        pixel_data[46][33] = 13;
        pixel_data[46][34] = 13;
        pixel_data[46][35] = 13;
        pixel_data[46][36] = 13;
        pixel_data[46][37] = 13;
        pixel_data[46][38] = 13;
        pixel_data[46][39] = 13;
        pixel_data[46][40] = 13;
        pixel_data[46][41] = 13;
        pixel_data[46][42] = 13;
        pixel_data[46][43] = 13;
        pixel_data[46][44] = 13;
        pixel_data[46][45] = 7;
        pixel_data[46][46] = 12;
        pixel_data[46][47] = 0;
        pixel_data[46][48] = 0;
        pixel_data[46][49] = 0; // y=46
        pixel_data[47][0] = 0;
        pixel_data[47][1] = 0;
        pixel_data[47][2] = 0;
        pixel_data[47][3] = 0;
        pixel_data[47][4] = 14;
        pixel_data[47][5] = 14;
        pixel_data[47][6] = 0;
        pixel_data[47][7] = 0;
        pixel_data[47][8] = 0;
        pixel_data[47][9] = 0;
        pixel_data[47][10] = 14;
        pixel_data[47][11] = 14;
        pixel_data[47][12] = 10;
        pixel_data[47][13] = 15;
        pixel_data[47][14] = 13;
        pixel_data[47][15] = 12;
        pixel_data[47][16] = 3;
        pixel_data[47][17] = 15;
        pixel_data[47][18] = 15;
        pixel_data[47][19] = 4;
        pixel_data[47][20] = 6;
        pixel_data[47][21] = 6;
        pixel_data[47][22] = 6;
        pixel_data[47][23] = 6;
        pixel_data[47][24] = 6;
        pixel_data[47][25] = 11;
        pixel_data[47][26] = 1;
        pixel_data[47][27] = 11;
        pixel_data[47][28] = 11;
        pixel_data[47][29] = 11;
        pixel_data[47][30] = 0;
        pixel_data[47][31] = 13;
        pixel_data[47][32] = 13;
        pixel_data[47][33] = 13;
        pixel_data[47][34] = 13;
        pixel_data[47][35] = 13;
        pixel_data[47][36] = 13;
        pixel_data[47][37] = 13;
        pixel_data[47][38] = 13;
        pixel_data[47][39] = 13;
        pixel_data[47][40] = 13;
        pixel_data[47][41] = 13;
        pixel_data[47][42] = 13;
        pixel_data[47][43] = 3;
        pixel_data[47][44] = 0;
        pixel_data[47][45] = 14;
        pixel_data[47][46] = 0;
        pixel_data[47][47] = 0;
        pixel_data[47][48] = 0;
        pixel_data[47][49] = 0; // y=47
        pixel_data[48][0] = 0;
        pixel_data[48][1] = 0;
        pixel_data[48][2] = 0;
        pixel_data[48][3] = 0;
        pixel_data[48][4] = 0;
        pixel_data[48][5] = 0;
        pixel_data[48][6] = 12;
        pixel_data[48][7] = 14;
        pixel_data[48][8] = 14;
        pixel_data[48][9] = 12;
        pixel_data[48][10] = 0;
        pixel_data[48][11] = 0;
        pixel_data[48][12] = 14;
        pixel_data[48][13] = 0;
        pixel_data[48][14] = 15;
        pixel_data[48][15] = 13;
        pixel_data[48][16] = 13;
        pixel_data[48][17] = 13;
        pixel_data[48][18] = 13;
        pixel_data[48][19] = 13;
        pixel_data[48][20] = 13;
        pixel_data[48][21] = 13;
        pixel_data[48][22] = 13;
        pixel_data[48][23] = 3;
        pixel_data[48][24] = 15;
        pixel_data[48][25] = 0;
        pixel_data[48][26] = 0;
        pixel_data[48][27] = 0;
        pixel_data[48][28] = 0;
        pixel_data[48][29] = 0;
        pixel_data[48][30] = 12;
        pixel_data[48][31] = 0;
        pixel_data[48][32] = 15;
        pixel_data[48][33] = 13;
        pixel_data[48][34] = 13;
        pixel_data[48][35] = 13;
        pixel_data[48][36] = 13;
        pixel_data[48][37] = 13;
        pixel_data[48][38] = 13;
        pixel_data[48][39] = 13;
        pixel_data[48][40] = 13;
        pixel_data[48][41] = 13;
        pixel_data[48][42] = 7;
        pixel_data[48][43] = 0;
        pixel_data[48][44] = 14;
        pixel_data[48][45] = 0;
        pixel_data[48][46] = 0;
        pixel_data[48][47] = 0;
        pixel_data[48][48] = 0;
        pixel_data[48][49] = 0; // y=48
        pixel_data[49][0] = 0;
        pixel_data[49][1] = 0;
        pixel_data[49][2] = 0;
        pixel_data[49][3] = 0;
        pixel_data[49][4] = 0;
        pixel_data[49][5] = 0;
        pixel_data[49][6] = 0;
        pixel_data[49][7] = 0;
        pixel_data[49][8] = 0;
        pixel_data[49][9] = 0;
        pixel_data[49][10] = 0;
        pixel_data[49][11] = 0;
        pixel_data[49][12] = 0;
        pixel_data[49][13] = 14;
        pixel_data[49][14] = 0;
        pixel_data[49][15] = 3;
        pixel_data[49][16] = 13;
        pixel_data[49][17] = 13;
        pixel_data[49][18] = 13;
        pixel_data[49][19] = 13;
        pixel_data[49][20] = 13;
        pixel_data[49][21] = 13;
        pixel_data[49][22] = 13;
        pixel_data[49][23] = 0;
        pixel_data[49][24] = 0;
        pixel_data[49][25] = 12;
        pixel_data[49][26] = 0;
        pixel_data[49][27] = 1;
        pixel_data[49][28] = 5;
        pixel_data[49][29] = 1;
        pixel_data[49][30] = 0;
        pixel_data[49][31] = 14;
        pixel_data[49][32] = 0;
        pixel_data[49][33] = 0;
        pixel_data[49][34] = 13;
        pixel_data[49][35] = 13;
        pixel_data[49][36] = 13;
        pixel_data[49][37] = 13;
        pixel_data[49][38] = 13;
        pixel_data[49][39] = 13;
        pixel_data[49][40] = 15;
        pixel_data[49][41] = 0;
        pixel_data[49][42] = 0;
        pixel_data[49][43] = 12;
        pixel_data[49][44] = 0;
        pixel_data[49][45] = 0;
        pixel_data[49][46] = 0;
        pixel_data[49][47] = 0;
        pixel_data[49][48] = 0;
        pixel_data[49][49] = 0; // y=49
    end
endmodule
