module bullet2_lut(output reg [3:0] pixel_data [0:99][0:99]);
    initial begin
        pixel_data[0][0] = 0;
        pixel_data[0][1] = 0;
        pixel_data[0][2] = 0;
        pixel_data[0][3] = 0;
        pixel_data[0][4] = 0;
        pixel_data[0][5] = 0;
        pixel_data[0][6] = 0;
        pixel_data[0][7] = 0;
        pixel_data[0][8] = 0;
        pixel_data[0][9] = 0;
        pixel_data[0][10] = 0;
        pixel_data[0][11] = 0;
        pixel_data[0][12] = 0;
        pixel_data[0][13] = 0;
        pixel_data[0][14] = 0;
        pixel_data[0][15] = 0;
        pixel_data[0][16] = 0;
        pixel_data[0][17] = 0;
        pixel_data[0][18] = 0;
        pixel_data[0][19] = 0;
        pixel_data[0][20] = 0;
        pixel_data[0][21] = 0;
        pixel_data[0][22] = 0;
        pixel_data[0][23] = 0;
        pixel_data[0][24] = 0;
        pixel_data[0][25] = 0;
        pixel_data[0][26] = 0;
        pixel_data[0][27] = 0;
        pixel_data[0][28] = 0;
        pixel_data[0][29] = 0;
        pixel_data[0][30] = 0;
        pixel_data[0][31] = 0;
        pixel_data[0][32] = 0;
        pixel_data[0][33] = 0;
        pixel_data[0][34] = 0;
        pixel_data[0][35] = 0;
        pixel_data[0][36] = 0;
        pixel_data[0][37] = 0;
        pixel_data[0][38] = 0;
        pixel_data[0][39] = 0;
        pixel_data[0][40] = 0;
        pixel_data[0][41] = 0;
        pixel_data[0][42] = 0;
        pixel_data[0][43] = 0;
        pixel_data[0][44] = 0;
        pixel_data[0][45] = 0;
        pixel_data[0][46] = 0;
        pixel_data[0][47] = 0;
        pixel_data[0][48] = 0;
        pixel_data[0][49] = 0;
        pixel_data[0][50] = 0;
        pixel_data[0][51] = 0;
        pixel_data[0][52] = 0;
        pixel_data[0][53] = 0;
        pixel_data[0][54] = 0;
        pixel_data[0][55] = 0;
        pixel_data[0][56] = 0;
        pixel_data[0][57] = 0;
        pixel_data[0][58] = 0;
        pixel_data[0][59] = 0;
        pixel_data[0][60] = 0;
        pixel_data[0][61] = 0;
        pixel_data[0][62] = 0;
        pixel_data[0][63] = 0;
        pixel_data[0][64] = 0;
        pixel_data[0][65] = 0;
        pixel_data[0][66] = 0;
        pixel_data[0][67] = 0;
        pixel_data[0][68] = 0;
        pixel_data[0][69] = 0;
        pixel_data[0][70] = 0;
        pixel_data[0][71] = 0;
        pixel_data[0][72] = 0;
        pixel_data[0][73] = 0;
        pixel_data[0][74] = 0;
        pixel_data[0][75] = 0;
        pixel_data[0][76] = 0;
        pixel_data[0][77] = 0;
        pixel_data[0][78] = 0;
        pixel_data[0][79] = 0;
        pixel_data[0][80] = 0;
        pixel_data[0][81] = 0;
        pixel_data[0][82] = 0;
        pixel_data[0][83] = 0;
        pixel_data[0][84] = 0;
        pixel_data[0][85] = 0;
        pixel_data[0][86] = 0;
        pixel_data[0][87] = 0;
        pixel_data[0][88] = 0;
        pixel_data[0][89] = 0;
        pixel_data[0][90] = 0;
        pixel_data[0][91] = 0;
        pixel_data[0][92] = 0;
        pixel_data[0][93] = 0;
        pixel_data[0][94] = 0;
        pixel_data[0][95] = 0;
        pixel_data[0][96] = 0;
        pixel_data[0][97] = 0;
        pixel_data[0][98] = 0;
        pixel_data[0][99] = 0; // y=0
        pixel_data[1][0] = 0;
        pixel_data[1][1] = 0;
        pixel_data[1][2] = 0;
        pixel_data[1][3] = 0;
        pixel_data[1][4] = 0;
        pixel_data[1][5] = 0;
        pixel_data[1][6] = 0;
        pixel_data[1][7] = 0;
        pixel_data[1][8] = 0;
        pixel_data[1][9] = 0;
        pixel_data[1][10] = 0;
        pixel_data[1][11] = 0;
        pixel_data[1][12] = 0;
        pixel_data[1][13] = 0;
        pixel_data[1][14] = 0;
        pixel_data[1][15] = 0;
        pixel_data[1][16] = 0;
        pixel_data[1][17] = 0;
        pixel_data[1][18] = 0;
        pixel_data[1][19] = 0;
        pixel_data[1][20] = 0;
        pixel_data[1][21] = 0;
        pixel_data[1][22] = 0;
        pixel_data[1][23] = 0;
        pixel_data[1][24] = 0;
        pixel_data[1][25] = 0;
        pixel_data[1][26] = 0;
        pixel_data[1][27] = 0;
        pixel_data[1][28] = 0;
        pixel_data[1][29] = 0;
        pixel_data[1][30] = 0;
        pixel_data[1][31] = 0;
        pixel_data[1][32] = 0;
        pixel_data[1][33] = 0;
        pixel_data[1][34] = 0;
        pixel_data[1][35] = 0;
        pixel_data[1][36] = 0;
        pixel_data[1][37] = 0;
        pixel_data[1][38] = 0;
        pixel_data[1][39] = 0;
        pixel_data[1][40] = 0;
        pixel_data[1][41] = 0;
        pixel_data[1][42] = 0;
        pixel_data[1][43] = 0;
        pixel_data[1][44] = 0;
        pixel_data[1][45] = 0;
        pixel_data[1][46] = 0;
        pixel_data[1][47] = 0;
        pixel_data[1][48] = 0;
        pixel_data[1][49] = 0;
        pixel_data[1][50] = 0;
        pixel_data[1][51] = 0;
        pixel_data[1][52] = 0;
        pixel_data[1][53] = 0;
        pixel_data[1][54] = 0;
        pixel_data[1][55] = 0;
        pixel_data[1][56] = 0;
        pixel_data[1][57] = 0;
        pixel_data[1][58] = 0;
        pixel_data[1][59] = 0;
        pixel_data[1][60] = 0;
        pixel_data[1][61] = 0;
        pixel_data[1][62] = 0;
        pixel_data[1][63] = 0;
        pixel_data[1][64] = 0;
        pixel_data[1][65] = 0;
        pixel_data[1][66] = 0;
        pixel_data[1][67] = 0;
        pixel_data[1][68] = 0;
        pixel_data[1][69] = 0;
        pixel_data[1][70] = 0;
        pixel_data[1][71] = 0;
        pixel_data[1][72] = 0;
        pixel_data[1][73] = 0;
        pixel_data[1][74] = 0;
        pixel_data[1][75] = 0;
        pixel_data[1][76] = 0;
        pixel_data[1][77] = 0;
        pixel_data[1][78] = 0;
        pixel_data[1][79] = 0;
        pixel_data[1][80] = 0;
        pixel_data[1][81] = 0;
        pixel_data[1][82] = 0;
        pixel_data[1][83] = 0;
        pixel_data[1][84] = 0;
        pixel_data[1][85] = 0;
        pixel_data[1][86] = 0;
        pixel_data[1][87] = 0;
        pixel_data[1][88] = 0;
        pixel_data[1][89] = 0;
        pixel_data[1][90] = 0;
        pixel_data[1][91] = 0;
        pixel_data[1][92] = 0;
        pixel_data[1][93] = 0;
        pixel_data[1][94] = 0;
        pixel_data[1][95] = 0;
        pixel_data[1][96] = 0;
        pixel_data[1][97] = 0;
        pixel_data[1][98] = 0;
        pixel_data[1][99] = 0; // y=1
        pixel_data[2][0] = 0;
        pixel_data[2][1] = 0;
        pixel_data[2][2] = 0;
        pixel_data[2][3] = 0;
        pixel_data[2][4] = 0;
        pixel_data[2][5] = 0;
        pixel_data[2][6] = 0;
        pixel_data[2][7] = 0;
        pixel_data[2][8] = 0;
        pixel_data[2][9] = 0;
        pixel_data[2][10] = 0;
        pixel_data[2][11] = 0;
        pixel_data[2][12] = 0;
        pixel_data[2][13] = 0;
        pixel_data[2][14] = 0;
        pixel_data[2][15] = 0;
        pixel_data[2][16] = 0;
        pixel_data[2][17] = 0;
        pixel_data[2][18] = 0;
        pixel_data[2][19] = 0;
        pixel_data[2][20] = 0;
        pixel_data[2][21] = 0;
        pixel_data[2][22] = 0;
        pixel_data[2][23] = 0;
        pixel_data[2][24] = 0;
        pixel_data[2][25] = 0;
        pixel_data[2][26] = 0;
        pixel_data[2][27] = 0;
        pixel_data[2][28] = 0;
        pixel_data[2][29] = 0;
        pixel_data[2][30] = 0;
        pixel_data[2][31] = 0;
        pixel_data[2][32] = 0;
        pixel_data[2][33] = 0;
        pixel_data[2][34] = 0;
        pixel_data[2][35] = 0;
        pixel_data[2][36] = 0;
        pixel_data[2][37] = 0;
        pixel_data[2][38] = 0;
        pixel_data[2][39] = 0;
        pixel_data[2][40] = 0;
        pixel_data[2][41] = 0;
        pixel_data[2][42] = 0;
        pixel_data[2][43] = 0;
        pixel_data[2][44] = 0;
        pixel_data[2][45] = 0;
        pixel_data[2][46] = 0;
        pixel_data[2][47] = 0;
        pixel_data[2][48] = 0;
        pixel_data[2][49] = 0;
        pixel_data[2][50] = 0;
        pixel_data[2][51] = 0;
        pixel_data[2][52] = 0;
        pixel_data[2][53] = 0;
        pixel_data[2][54] = 0;
        pixel_data[2][55] = 0;
        pixel_data[2][56] = 0;
        pixel_data[2][57] = 0;
        pixel_data[2][58] = 0;
        pixel_data[2][59] = 0;
        pixel_data[2][60] = 0;
        pixel_data[2][61] = 0;
        pixel_data[2][62] = 0;
        pixel_data[2][63] = 0;
        pixel_data[2][64] = 0;
        pixel_data[2][65] = 0;
        pixel_data[2][66] = 0;
        pixel_data[2][67] = 0;
        pixel_data[2][68] = 0;
        pixel_data[2][69] = 0;
        pixel_data[2][70] = 0;
        pixel_data[2][71] = 0;
        pixel_data[2][72] = 0;
        pixel_data[2][73] = 0;
        pixel_data[2][74] = 0;
        pixel_data[2][75] = 0;
        pixel_data[2][76] = 0;
        pixel_data[2][77] = 0;
        pixel_data[2][78] = 0;
        pixel_data[2][79] = 0;
        pixel_data[2][80] = 0;
        pixel_data[2][81] = 0;
        pixel_data[2][82] = 0;
        pixel_data[2][83] = 0;
        pixel_data[2][84] = 0;
        pixel_data[2][85] = 0;
        pixel_data[2][86] = 0;
        pixel_data[2][87] = 0;
        pixel_data[2][88] = 0;
        pixel_data[2][89] = 0;
        pixel_data[2][90] = 0;
        pixel_data[2][91] = 0;
        pixel_data[2][92] = 0;
        pixel_data[2][93] = 0;
        pixel_data[2][94] = 0;
        pixel_data[2][95] = 0;
        pixel_data[2][96] = 0;
        pixel_data[2][97] = 0;
        pixel_data[2][98] = 0;
        pixel_data[2][99] = 0; // y=2
        pixel_data[3][0] = 0;
        pixel_data[3][1] = 0;
        pixel_data[3][2] = 0;
        pixel_data[3][3] = 0;
        pixel_data[3][4] = 0;
        pixel_data[3][5] = 0;
        pixel_data[3][6] = 0;
        pixel_data[3][7] = 0;
        pixel_data[3][8] = 0;
        pixel_data[3][9] = 0;
        pixel_data[3][10] = 0;
        pixel_data[3][11] = 0;
        pixel_data[3][12] = 0;
        pixel_data[3][13] = 0;
        pixel_data[3][14] = 0;
        pixel_data[3][15] = 0;
        pixel_data[3][16] = 0;
        pixel_data[3][17] = 0;
        pixel_data[3][18] = 0;
        pixel_data[3][19] = 0;
        pixel_data[3][20] = 0;
        pixel_data[3][21] = 0;
        pixel_data[3][22] = 0;
        pixel_data[3][23] = 0;
        pixel_data[3][24] = 0;
        pixel_data[3][25] = 0;
        pixel_data[3][26] = 0;
        pixel_data[3][27] = 0;
        pixel_data[3][28] = 0;
        pixel_data[3][29] = 0;
        pixel_data[3][30] = 0;
        pixel_data[3][31] = 0;
        pixel_data[3][32] = 0;
        pixel_data[3][33] = 0;
        pixel_data[3][34] = 0;
        pixel_data[3][35] = 0;
        pixel_data[3][36] = 0;
        pixel_data[3][37] = 0;
        pixel_data[3][38] = 0;
        pixel_data[3][39] = 0;
        pixel_data[3][40] = 0;
        pixel_data[3][41] = 0;
        pixel_data[3][42] = 0;
        pixel_data[3][43] = 0;
        pixel_data[3][44] = 0;
        pixel_data[3][45] = 0;
        pixel_data[3][46] = 0;
        pixel_data[3][47] = 0;
        pixel_data[3][48] = 0;
        pixel_data[3][49] = 0;
        pixel_data[3][50] = 0;
        pixel_data[3][51] = 0;
        pixel_data[3][52] = 0;
        pixel_data[3][53] = 0;
        pixel_data[3][54] = 0;
        pixel_data[3][55] = 0;
        pixel_data[3][56] = 0;
        pixel_data[3][57] = 0;
        pixel_data[3][58] = 0;
        pixel_data[3][59] = 0;
        pixel_data[3][60] = 0;
        pixel_data[3][61] = 0;
        pixel_data[3][62] = 0;
        pixel_data[3][63] = 0;
        pixel_data[3][64] = 0;
        pixel_data[3][65] = 0;
        pixel_data[3][66] = 0;
        pixel_data[3][67] = 0;
        pixel_data[3][68] = 0;
        pixel_data[3][69] = 0;
        pixel_data[3][70] = 0;
        pixel_data[3][71] = 0;
        pixel_data[3][72] = 0;
        pixel_data[3][73] = 0;
        pixel_data[3][74] = 0;
        pixel_data[3][75] = 0;
        pixel_data[3][76] = 0;
        pixel_data[3][77] = 0;
        pixel_data[3][78] = 0;
        pixel_data[3][79] = 0;
        pixel_data[3][80] = 0;
        pixel_data[3][81] = 0;
        pixel_data[3][82] = 0;
        pixel_data[3][83] = 0;
        pixel_data[3][84] = 0;
        pixel_data[3][85] = 0;
        pixel_data[3][86] = 0;
        pixel_data[3][87] = 0;
        pixel_data[3][88] = 0;
        pixel_data[3][89] = 0;
        pixel_data[3][90] = 0;
        pixel_data[3][91] = 0;
        pixel_data[3][92] = 0;
        pixel_data[3][93] = 0;
        pixel_data[3][94] = 0;
        pixel_data[3][95] = 0;
        pixel_data[3][96] = 0;
        pixel_data[3][97] = 0;
        pixel_data[3][98] = 0;
        pixel_data[3][99] = 0; // y=3
        pixel_data[4][0] = 0;
        pixel_data[4][1] = 0;
        pixel_data[4][2] = 0;
        pixel_data[4][3] = 0;
        pixel_data[4][4] = 0;
        pixel_data[4][5] = 0;
        pixel_data[4][6] = 0;
        pixel_data[4][7] = 0;
        pixel_data[4][8] = 0;
        pixel_data[4][9] = 0;
        pixel_data[4][10] = 0;
        pixel_data[4][11] = 0;
        pixel_data[4][12] = 0;
        pixel_data[4][13] = 0;
        pixel_data[4][14] = 0;
        pixel_data[4][15] = 0;
        pixel_data[4][16] = 0;
        pixel_data[4][17] = 0;
        pixel_data[4][18] = 0;
        pixel_data[4][19] = 0;
        pixel_data[4][20] = 0;
        pixel_data[4][21] = 0;
        pixel_data[4][22] = 0;
        pixel_data[4][23] = 0;
        pixel_data[4][24] = 0;
        pixel_data[4][25] = 0;
        pixel_data[4][26] = 0;
        pixel_data[4][27] = 0;
        pixel_data[4][28] = 0;
        pixel_data[4][29] = 0;
        pixel_data[4][30] = 0;
        pixel_data[4][31] = 0;
        pixel_data[4][32] = 0;
        pixel_data[4][33] = 0;
        pixel_data[4][34] = 0;
        pixel_data[4][35] = 0;
        pixel_data[4][36] = 0;
        pixel_data[4][37] = 0;
        pixel_data[4][38] = 0;
        pixel_data[4][39] = 0;
        pixel_data[4][40] = 0;
        pixel_data[4][41] = 0;
        pixel_data[4][42] = 0;
        pixel_data[4][43] = 0;
        pixel_data[4][44] = 0;
        pixel_data[4][45] = 0;
        pixel_data[4][46] = 0;
        pixel_data[4][47] = 0;
        pixel_data[4][48] = 0;
        pixel_data[4][49] = 0;
        pixel_data[4][50] = 0;
        pixel_data[4][51] = 0;
        pixel_data[4][52] = 0;
        pixel_data[4][53] = 0;
        pixel_data[4][54] = 0;
        pixel_data[4][55] = 0;
        pixel_data[4][56] = 0;
        pixel_data[4][57] = 0;
        pixel_data[4][58] = 0;
        pixel_data[4][59] = 0;
        pixel_data[4][60] = 0;
        pixel_data[4][61] = 0;
        pixel_data[4][62] = 0;
        pixel_data[4][63] = 0;
        pixel_data[4][64] = 0;
        pixel_data[4][65] = 0;
        pixel_data[4][66] = 0;
        pixel_data[4][67] = 0;
        pixel_data[4][68] = 0;
        pixel_data[4][69] = 0;
        pixel_data[4][70] = 0;
        pixel_data[4][71] = 0;
        pixel_data[4][72] = 0;
        pixel_data[4][73] = 0;
        pixel_data[4][74] = 0;
        pixel_data[4][75] = 0;
        pixel_data[4][76] = 0;
        pixel_data[4][77] = 0;
        pixel_data[4][78] = 0;
        pixel_data[4][79] = 0;
        pixel_data[4][80] = 0;
        pixel_data[4][81] = 0;
        pixel_data[4][82] = 0;
        pixel_data[4][83] = 0;
        pixel_data[4][84] = 0;
        pixel_data[4][85] = 0;
        pixel_data[4][86] = 0;
        pixel_data[4][87] = 0;
        pixel_data[4][88] = 0;
        pixel_data[4][89] = 0;
        pixel_data[4][90] = 0;
        pixel_data[4][91] = 0;
        pixel_data[4][92] = 0;
        pixel_data[4][93] = 0;
        pixel_data[4][94] = 0;
        pixel_data[4][95] = 0;
        pixel_data[4][96] = 0;
        pixel_data[4][97] = 0;
        pixel_data[4][98] = 0;
        pixel_data[4][99] = 0; // y=4
        pixel_data[5][0] = 0;
        pixel_data[5][1] = 0;
        pixel_data[5][2] = 0;
        pixel_data[5][3] = 0;
        pixel_data[5][4] = 0;
        pixel_data[5][5] = 0;
        pixel_data[5][6] = 0;
        pixel_data[5][7] = 0;
        pixel_data[5][8] = 0;
        pixel_data[5][9] = 0;
        pixel_data[5][10] = 0;
        pixel_data[5][11] = 0;
        pixel_data[5][12] = 0;
        pixel_data[5][13] = 0;
        pixel_data[5][14] = 0;
        pixel_data[5][15] = 0;
        pixel_data[5][16] = 0;
        pixel_data[5][17] = 0;
        pixel_data[5][18] = 0;
        pixel_data[5][19] = 0;
        pixel_data[5][20] = 0;
        pixel_data[5][21] = 0;
        pixel_data[5][22] = 0;
        pixel_data[5][23] = 0;
        pixel_data[5][24] = 0;
        pixel_data[5][25] = 0;
        pixel_data[5][26] = 0;
        pixel_data[5][27] = 0;
        pixel_data[5][28] = 0;
        pixel_data[5][29] = 0;
        pixel_data[5][30] = 0;
        pixel_data[5][31] = 0;
        pixel_data[5][32] = 0;
        pixel_data[5][33] = 0;
        pixel_data[5][34] = 0;
        pixel_data[5][35] = 0;
        pixel_data[5][36] = 0;
        pixel_data[5][37] = 0;
        pixel_data[5][38] = 0;
        pixel_data[5][39] = 0;
        pixel_data[5][40] = 0;
        pixel_data[5][41] = 0;
        pixel_data[5][42] = 0;
        pixel_data[5][43] = 0;
        pixel_data[5][44] = 0;
        pixel_data[5][45] = 0;
        pixel_data[5][46] = 0;
        pixel_data[5][47] = 0;
        pixel_data[5][48] = 0;
        pixel_data[5][49] = 0;
        pixel_data[5][50] = 0;
        pixel_data[5][51] = 0;
        pixel_data[5][52] = 0;
        pixel_data[5][53] = 0;
        pixel_data[5][54] = 0;
        pixel_data[5][55] = 0;
        pixel_data[5][56] = 0;
        pixel_data[5][57] = 0;
        pixel_data[5][58] = 0;
        pixel_data[5][59] = 0;
        pixel_data[5][60] = 0;
        pixel_data[5][61] = 0;
        pixel_data[5][62] = 0;
        pixel_data[5][63] = 0;
        pixel_data[5][64] = 0;
        pixel_data[5][65] = 0;
        pixel_data[5][66] = 0;
        pixel_data[5][67] = 0;
        pixel_data[5][68] = 0;
        pixel_data[5][69] = 0;
        pixel_data[5][70] = 0;
        pixel_data[5][71] = 0;
        pixel_data[5][72] = 0;
        pixel_data[5][73] = 0;
        pixel_data[5][74] = 0;
        pixel_data[5][75] = 0;
        pixel_data[5][76] = 0;
        pixel_data[5][77] = 0;
        pixel_data[5][78] = 0;
        pixel_data[5][79] = 0;
        pixel_data[5][80] = 0;
        pixel_data[5][81] = 0;
        pixel_data[5][82] = 0;
        pixel_data[5][83] = 0;
        pixel_data[5][84] = 0;
        pixel_data[5][85] = 0;
        pixel_data[5][86] = 0;
        pixel_data[5][87] = 0;
        pixel_data[5][88] = 0;
        pixel_data[5][89] = 0;
        pixel_data[5][90] = 0;
        pixel_data[5][91] = 0;
        pixel_data[5][92] = 0;
        pixel_data[5][93] = 0;
        pixel_data[5][94] = 0;
        pixel_data[5][95] = 0;
        pixel_data[5][96] = 0;
        pixel_data[5][97] = 0;
        pixel_data[5][98] = 0;
        pixel_data[5][99] = 0; // y=5
        pixel_data[6][0] = 0;
        pixel_data[6][1] = 0;
        pixel_data[6][2] = 0;
        pixel_data[6][3] = 0;
        pixel_data[6][4] = 0;
        pixel_data[6][5] = 0;
        pixel_data[6][6] = 0;
        pixel_data[6][7] = 0;
        pixel_data[6][8] = 0;
        pixel_data[6][9] = 0;
        pixel_data[6][10] = 0;
        pixel_data[6][11] = 0;
        pixel_data[6][12] = 0;
        pixel_data[6][13] = 0;
        pixel_data[6][14] = 0;
        pixel_data[6][15] = 0;
        pixel_data[6][16] = 0;
        pixel_data[6][17] = 0;
        pixel_data[6][18] = 0;
        pixel_data[6][19] = 0;
        pixel_data[6][20] = 0;
        pixel_data[6][21] = 0;
        pixel_data[6][22] = 0;
        pixel_data[6][23] = 0;
        pixel_data[6][24] = 0;
        pixel_data[6][25] = 0;
        pixel_data[6][26] = 0;
        pixel_data[6][27] = 0;
        pixel_data[6][28] = 0;
        pixel_data[6][29] = 0;
        pixel_data[6][30] = 0;
        pixel_data[6][31] = 0;
        pixel_data[6][32] = 0;
        pixel_data[6][33] = 0;
        pixel_data[6][34] = 0;
        pixel_data[6][35] = 0;
        pixel_data[6][36] = 0;
        pixel_data[6][37] = 0;
        pixel_data[6][38] = 0;
        pixel_data[6][39] = 0;
        pixel_data[6][40] = 0;
        pixel_data[6][41] = 0;
        pixel_data[6][42] = 0;
        pixel_data[6][43] = 0;
        pixel_data[6][44] = 0;
        pixel_data[6][45] = 0;
        pixel_data[6][46] = 0;
        pixel_data[6][47] = 0;
        pixel_data[6][48] = 0;
        pixel_data[6][49] = 0;
        pixel_data[6][50] = 0;
        pixel_data[6][51] = 0;
        pixel_data[6][52] = 0;
        pixel_data[6][53] = 0;
        pixel_data[6][54] = 0;
        pixel_data[6][55] = 0;
        pixel_data[6][56] = 0;
        pixel_data[6][57] = 0;
        pixel_data[6][58] = 0;
        pixel_data[6][59] = 0;
        pixel_data[6][60] = 0;
        pixel_data[6][61] = 0;
        pixel_data[6][62] = 0;
        pixel_data[6][63] = 0;
        pixel_data[6][64] = 0;
        pixel_data[6][65] = 0;
        pixel_data[6][66] = 0;
        pixel_data[6][67] = 0;
        pixel_data[6][68] = 0;
        pixel_data[6][69] = 0;
        pixel_data[6][70] = 0;
        pixel_data[6][71] = 0;
        pixel_data[6][72] = 0;
        pixel_data[6][73] = 0;
        pixel_data[6][74] = 0;
        pixel_data[6][75] = 0;
        pixel_data[6][76] = 0;
        pixel_data[6][77] = 0;
        pixel_data[6][78] = 0;
        pixel_data[6][79] = 0;
        pixel_data[6][80] = 0;
        pixel_data[6][81] = 0;
        pixel_data[6][82] = 0;
        pixel_data[6][83] = 0;
        pixel_data[6][84] = 0;
        pixel_data[6][85] = 0;
        pixel_data[6][86] = 0;
        pixel_data[6][87] = 0;
        pixel_data[6][88] = 0;
        pixel_data[6][89] = 0;
        pixel_data[6][90] = 0;
        pixel_data[6][91] = 0;
        pixel_data[6][92] = 0;
        pixel_data[6][93] = 0;
        pixel_data[6][94] = 0;
        pixel_data[6][95] = 0;
        pixel_data[6][96] = 0;
        pixel_data[6][97] = 0;
        pixel_data[6][98] = 0;
        pixel_data[6][99] = 0; // y=6
        pixel_data[7][0] = 0;
        pixel_data[7][1] = 0;
        pixel_data[7][2] = 0;
        pixel_data[7][3] = 0;
        pixel_data[7][4] = 0;
        pixel_data[7][5] = 0;
        pixel_data[7][6] = 0;
        pixel_data[7][7] = 0;
        pixel_data[7][8] = 0;
        pixel_data[7][9] = 0;
        pixel_data[7][10] = 0;
        pixel_data[7][11] = 0;
        pixel_data[7][12] = 0;
        pixel_data[7][13] = 0;
        pixel_data[7][14] = 0;
        pixel_data[7][15] = 0;
        pixel_data[7][16] = 0;
        pixel_data[7][17] = 0;
        pixel_data[7][18] = 0;
        pixel_data[7][19] = 0;
        pixel_data[7][20] = 0;
        pixel_data[7][21] = 0;
        pixel_data[7][22] = 0;
        pixel_data[7][23] = 0;
        pixel_data[7][24] = 0;
        pixel_data[7][25] = 0;
        pixel_data[7][26] = 0;
        pixel_data[7][27] = 0;
        pixel_data[7][28] = 0;
        pixel_data[7][29] = 0;
        pixel_data[7][30] = 0;
        pixel_data[7][31] = 0;
        pixel_data[7][32] = 0;
        pixel_data[7][33] = 0;
        pixel_data[7][34] = 0;
        pixel_data[7][35] = 0;
        pixel_data[7][36] = 0;
        pixel_data[7][37] = 0;
        pixel_data[7][38] = 0;
        pixel_data[7][39] = 0;
        pixel_data[7][40] = 0;
        pixel_data[7][41] = 0;
        pixel_data[7][42] = 0;
        pixel_data[7][43] = 0;
        pixel_data[7][44] = 0;
        pixel_data[7][45] = 0;
        pixel_data[7][46] = 0;
        pixel_data[7][47] = 0;
        pixel_data[7][48] = 0;
        pixel_data[7][49] = 0;
        pixel_data[7][50] = 0;
        pixel_data[7][51] = 0;
        pixel_data[7][52] = 0;
        pixel_data[7][53] = 0;
        pixel_data[7][54] = 0;
        pixel_data[7][55] = 0;
        pixel_data[7][56] = 0;
        pixel_data[7][57] = 0;
        pixel_data[7][58] = 0;
        pixel_data[7][59] = 0;
        pixel_data[7][60] = 0;
        pixel_data[7][61] = 0;
        pixel_data[7][62] = 0;
        pixel_data[7][63] = 0;
        pixel_data[7][64] = 0;
        pixel_data[7][65] = 0;
        pixel_data[7][66] = 0;
        pixel_data[7][67] = 0;
        pixel_data[7][68] = 0;
        pixel_data[7][69] = 0;
        pixel_data[7][70] = 0;
        pixel_data[7][71] = 0;
        pixel_data[7][72] = 0;
        pixel_data[7][73] = 0;
        pixel_data[7][74] = 0;
        pixel_data[7][75] = 0;
        pixel_data[7][76] = 0;
        pixel_data[7][77] = 0;
        pixel_data[7][78] = 0;
        pixel_data[7][79] = 0;
        pixel_data[7][80] = 0;
        pixel_data[7][81] = 0;
        pixel_data[7][82] = 0;
        pixel_data[7][83] = 0;
        pixel_data[7][84] = 0;
        pixel_data[7][85] = 0;
        pixel_data[7][86] = 0;
        pixel_data[7][87] = 0;
        pixel_data[7][88] = 0;
        pixel_data[7][89] = 0;
        pixel_data[7][90] = 0;
        pixel_data[7][91] = 0;
        pixel_data[7][92] = 0;
        pixel_data[7][93] = 0;
        pixel_data[7][94] = 0;
        pixel_data[7][95] = 0;
        pixel_data[7][96] = 0;
        pixel_data[7][97] = 0;
        pixel_data[7][98] = 0;
        pixel_data[7][99] = 0; // y=7
        pixel_data[8][0] = 0;
        pixel_data[8][1] = 0;
        pixel_data[8][2] = 0;
        pixel_data[8][3] = 0;
        pixel_data[8][4] = 0;
        pixel_data[8][5] = 0;
        pixel_data[8][6] = 0;
        pixel_data[8][7] = 0;
        pixel_data[8][8] = 0;
        pixel_data[8][9] = 0;
        pixel_data[8][10] = 0;
        pixel_data[8][11] = 0;
        pixel_data[8][12] = 0;
        pixel_data[8][13] = 0;
        pixel_data[8][14] = 0;
        pixel_data[8][15] = 0;
        pixel_data[8][16] = 0;
        pixel_data[8][17] = 0;
        pixel_data[8][18] = 0;
        pixel_data[8][19] = 0;
        pixel_data[8][20] = 0;
        pixel_data[8][21] = 0;
        pixel_data[8][22] = 0;
        pixel_data[8][23] = 0;
        pixel_data[8][24] = 0;
        pixel_data[8][25] = 0;
        pixel_data[8][26] = 0;
        pixel_data[8][27] = 0;
        pixel_data[8][28] = 0;
        pixel_data[8][29] = 0;
        pixel_data[8][30] = 0;
        pixel_data[8][31] = 0;
        pixel_data[8][32] = 0;
        pixel_data[8][33] = 0;
        pixel_data[8][34] = 0;
        pixel_data[8][35] = 0;
        pixel_data[8][36] = 0;
        pixel_data[8][37] = 0;
        pixel_data[8][38] = 0;
        pixel_data[8][39] = 0;
        pixel_data[8][40] = 0;
        pixel_data[8][41] = 0;
        pixel_data[8][42] = 0;
        pixel_data[8][43] = 0;
        pixel_data[8][44] = 0;
        pixel_data[8][45] = 0;
        pixel_data[8][46] = 0;
        pixel_data[8][47] = 0;
        pixel_data[8][48] = 0;
        pixel_data[8][49] = 0;
        pixel_data[8][50] = 0;
        pixel_data[8][51] = 0;
        pixel_data[8][52] = 0;
        pixel_data[8][53] = 0;
        pixel_data[8][54] = 0;
        pixel_data[8][55] = 0;
        pixel_data[8][56] = 0;
        pixel_data[8][57] = 0;
        pixel_data[8][58] = 0;
        pixel_data[8][59] = 0;
        pixel_data[8][60] = 0;
        pixel_data[8][61] = 0;
        pixel_data[8][62] = 0;
        pixel_data[8][63] = 0;
        pixel_data[8][64] = 0;
        pixel_data[8][65] = 0;
        pixel_data[8][66] = 0;
        pixel_data[8][67] = 0;
        pixel_data[8][68] = 0;
        pixel_data[8][69] = 0;
        pixel_data[8][70] = 0;
        pixel_data[8][71] = 0;
        pixel_data[8][72] = 0;
        pixel_data[8][73] = 0;
        pixel_data[8][74] = 0;
        pixel_data[8][75] = 0;
        pixel_data[8][76] = 0;
        pixel_data[8][77] = 0;
        pixel_data[8][78] = 0;
        pixel_data[8][79] = 0;
        pixel_data[8][80] = 0;
        pixel_data[8][81] = 0;
        pixel_data[8][82] = 0;
        pixel_data[8][83] = 0;
        pixel_data[8][84] = 0;
        pixel_data[8][85] = 0;
        pixel_data[8][86] = 0;
        pixel_data[8][87] = 0;
        pixel_data[8][88] = 0;
        pixel_data[8][89] = 0;
        pixel_data[8][90] = 0;
        pixel_data[8][91] = 0;
        pixel_data[8][92] = 0;
        pixel_data[8][93] = 0;
        pixel_data[8][94] = 0;
        pixel_data[8][95] = 0;
        pixel_data[8][96] = 0;
        pixel_data[8][97] = 0;
        pixel_data[8][98] = 0;
        pixel_data[8][99] = 0; // y=8
        pixel_data[9][0] = 0;
        pixel_data[9][1] = 0;
        pixel_data[9][2] = 0;
        pixel_data[9][3] = 0;
        pixel_data[9][4] = 0;
        pixel_data[9][5] = 0;
        pixel_data[9][6] = 0;
        pixel_data[9][7] = 0;
        pixel_data[9][8] = 0;
        pixel_data[9][9] = 0;
        pixel_data[9][10] = 0;
        pixel_data[9][11] = 0;
        pixel_data[9][12] = 0;
        pixel_data[9][13] = 0;
        pixel_data[9][14] = 0;
        pixel_data[9][15] = 0;
        pixel_data[9][16] = 0;
        pixel_data[9][17] = 0;
        pixel_data[9][18] = 0;
        pixel_data[9][19] = 0;
        pixel_data[9][20] = 0;
        pixel_data[9][21] = 0;
        pixel_data[9][22] = 0;
        pixel_data[9][23] = 0;
        pixel_data[9][24] = 0;
        pixel_data[9][25] = 0;
        pixel_data[9][26] = 0;
        pixel_data[9][27] = 0;
        pixel_data[9][28] = 0;
        pixel_data[9][29] = 0;
        pixel_data[9][30] = 0;
        pixel_data[9][31] = 0;
        pixel_data[9][32] = 0;
        pixel_data[9][33] = 0;
        pixel_data[9][34] = 0;
        pixel_data[9][35] = 0;
        pixel_data[9][36] = 0;
        pixel_data[9][37] = 0;
        pixel_data[9][38] = 0;
        pixel_data[9][39] = 0;
        pixel_data[9][40] = 0;
        pixel_data[9][41] = 0;
        pixel_data[9][42] = 0;
        pixel_data[9][43] = 0;
        pixel_data[9][44] = 0;
        pixel_data[9][45] = 0;
        pixel_data[9][46] = 0;
        pixel_data[9][47] = 0;
        pixel_data[9][48] = 0;
        pixel_data[9][49] = 0;
        pixel_data[9][50] = 0;
        pixel_data[9][51] = 0;
        pixel_data[9][52] = 0;
        pixel_data[9][53] = 0;
        pixel_data[9][54] = 0;
        pixel_data[9][55] = 0;
        pixel_data[9][56] = 0;
        pixel_data[9][57] = 0;
        pixel_data[9][58] = 0;
        pixel_data[9][59] = 0;
        pixel_data[9][60] = 0;
        pixel_data[9][61] = 0;
        pixel_data[9][62] = 0;
        pixel_data[9][63] = 0;
        pixel_data[9][64] = 0;
        pixel_data[9][65] = 0;
        pixel_data[9][66] = 0;
        pixel_data[9][67] = 0;
        pixel_data[9][68] = 0;
        pixel_data[9][69] = 0;
        pixel_data[9][70] = 0;
        pixel_data[9][71] = 0;
        pixel_data[9][72] = 0;
        pixel_data[9][73] = 0;
        pixel_data[9][74] = 0;
        pixel_data[9][75] = 0;
        pixel_data[9][76] = 0;
        pixel_data[9][77] = 0;
        pixel_data[9][78] = 0;
        pixel_data[9][79] = 0;
        pixel_data[9][80] = 0;
        pixel_data[9][81] = 0;
        pixel_data[9][82] = 0;
        pixel_data[9][83] = 0;
        pixel_data[9][84] = 0;
        pixel_data[9][85] = 0;
        pixel_data[9][86] = 0;
        pixel_data[9][87] = 0;
        pixel_data[9][88] = 0;
        pixel_data[9][89] = 0;
        pixel_data[9][90] = 0;
        pixel_data[9][91] = 0;
        pixel_data[9][92] = 0;
        pixel_data[9][93] = 0;
        pixel_data[9][94] = 0;
        pixel_data[9][95] = 0;
        pixel_data[9][96] = 0;
        pixel_data[9][97] = 0;
        pixel_data[9][98] = 0;
        pixel_data[9][99] = 0; // y=9
        pixel_data[10][0] = 0;
        pixel_data[10][1] = 0;
        pixel_data[10][2] = 0;
        pixel_data[10][3] = 0;
        pixel_data[10][4] = 0;
        pixel_data[10][5] = 0;
        pixel_data[10][6] = 0;
        pixel_data[10][7] = 0;
        pixel_data[10][8] = 0;
        pixel_data[10][9] = 0;
        pixel_data[10][10] = 0;
        pixel_data[10][11] = 0;
        pixel_data[10][12] = 0;
        pixel_data[10][13] = 0;
        pixel_data[10][14] = 0;
        pixel_data[10][15] = 0;
        pixel_data[10][16] = 0;
        pixel_data[10][17] = 0;
        pixel_data[10][18] = 0;
        pixel_data[10][19] = 0;
        pixel_data[10][20] = 0;
        pixel_data[10][21] = 0;
        pixel_data[10][22] = 0;
        pixel_data[10][23] = 0;
        pixel_data[10][24] = 0;
        pixel_data[10][25] = 0;
        pixel_data[10][26] = 0;
        pixel_data[10][27] = 0;
        pixel_data[10][28] = 0;
        pixel_data[10][29] = 0;
        pixel_data[10][30] = 0;
        pixel_data[10][31] = 0;
        pixel_data[10][32] = 0;
        pixel_data[10][33] = 0;
        pixel_data[10][34] = 0;
        pixel_data[10][35] = 0;
        pixel_data[10][36] = 0;
        pixel_data[10][37] = 0;
        pixel_data[10][38] = 0;
        pixel_data[10][39] = 0;
        pixel_data[10][40] = 0;
        pixel_data[10][41] = 0;
        pixel_data[10][42] = 0;
        pixel_data[10][43] = 0;
        pixel_data[10][44] = 0;
        pixel_data[10][45] = 0;
        pixel_data[10][46] = 0;
        pixel_data[10][47] = 0;
        pixel_data[10][48] = 0;
        pixel_data[10][49] = 0;
        pixel_data[10][50] = 0;
        pixel_data[10][51] = 0;
        pixel_data[10][52] = 0;
        pixel_data[10][53] = 0;
        pixel_data[10][54] = 0;
        pixel_data[10][55] = 0;
        pixel_data[10][56] = 0;
        pixel_data[10][57] = 0;
        pixel_data[10][58] = 0;
        pixel_data[10][59] = 0;
        pixel_data[10][60] = 0;
        pixel_data[10][61] = 0;
        pixel_data[10][62] = 0;
        pixel_data[10][63] = 0;
        pixel_data[10][64] = 0;
        pixel_data[10][65] = 0;
        pixel_data[10][66] = 0;
        pixel_data[10][67] = 0;
        pixel_data[10][68] = 0;
        pixel_data[10][69] = 0;
        pixel_data[10][70] = 0;
        pixel_data[10][71] = 0;
        pixel_data[10][72] = 0;
        pixel_data[10][73] = 0;
        pixel_data[10][74] = 0;
        pixel_data[10][75] = 0;
        pixel_data[10][76] = 0;
        pixel_data[10][77] = 0;
        pixel_data[10][78] = 0;
        pixel_data[10][79] = 0;
        pixel_data[10][80] = 0;
        pixel_data[10][81] = 0;
        pixel_data[10][82] = 0;
        pixel_data[10][83] = 0;
        pixel_data[10][84] = 0;
        pixel_data[10][85] = 0;
        pixel_data[10][86] = 0;
        pixel_data[10][87] = 0;
        pixel_data[10][88] = 0;
        pixel_data[10][89] = 0;
        pixel_data[10][90] = 0;
        pixel_data[10][91] = 0;
        pixel_data[10][92] = 0;
        pixel_data[10][93] = 0;
        pixel_data[10][94] = 0;
        pixel_data[10][95] = 0;
        pixel_data[10][96] = 0;
        pixel_data[10][97] = 0;
        pixel_data[10][98] = 0;
        pixel_data[10][99] = 0; // y=10
        pixel_data[11][0] = 0;
        pixel_data[11][1] = 0;
        pixel_data[11][2] = 0;
        pixel_data[11][3] = 0;
        pixel_data[11][4] = 0;
        pixel_data[11][5] = 0;
        pixel_data[11][6] = 0;
        pixel_data[11][7] = 0;
        pixel_data[11][8] = 0;
        pixel_data[11][9] = 0;
        pixel_data[11][10] = 0;
        pixel_data[11][11] = 0;
        pixel_data[11][12] = 0;
        pixel_data[11][13] = 0;
        pixel_data[11][14] = 0;
        pixel_data[11][15] = 0;
        pixel_data[11][16] = 0;
        pixel_data[11][17] = 0;
        pixel_data[11][18] = 0;
        pixel_data[11][19] = 0;
        pixel_data[11][20] = 0;
        pixel_data[11][21] = 0;
        pixel_data[11][22] = 0;
        pixel_data[11][23] = 0;
        pixel_data[11][24] = 0;
        pixel_data[11][25] = 0;
        pixel_data[11][26] = 0;
        pixel_data[11][27] = 0;
        pixel_data[11][28] = 0;
        pixel_data[11][29] = 0;
        pixel_data[11][30] = 0;
        pixel_data[11][31] = 0;
        pixel_data[11][32] = 0;
        pixel_data[11][33] = 0;
        pixel_data[11][34] = 0;
        pixel_data[11][35] = 0;
        pixel_data[11][36] = 0;
        pixel_data[11][37] = 0;
        pixel_data[11][38] = 0;
        pixel_data[11][39] = 0;
        pixel_data[11][40] = 0;
        pixel_data[11][41] = 0;
        pixel_data[11][42] = 0;
        pixel_data[11][43] = 0;
        pixel_data[11][44] = 0;
        pixel_data[11][45] = 0;
        pixel_data[11][46] = 0;
        pixel_data[11][47] = 0;
        pixel_data[11][48] = 0;
        pixel_data[11][49] = 0;
        pixel_data[11][50] = 0;
        pixel_data[11][51] = 0;
        pixel_data[11][52] = 0;
        pixel_data[11][53] = 0;
        pixel_data[11][54] = 0;
        pixel_data[11][55] = 0;
        pixel_data[11][56] = 0;
        pixel_data[11][57] = 0;
        pixel_data[11][58] = 0;
        pixel_data[11][59] = 0;
        pixel_data[11][60] = 0;
        pixel_data[11][61] = 0;
        pixel_data[11][62] = 0;
        pixel_data[11][63] = 0;
        pixel_data[11][64] = 0;
        pixel_data[11][65] = 0;
        pixel_data[11][66] = 0;
        pixel_data[11][67] = 0;
        pixel_data[11][68] = 0;
        pixel_data[11][69] = 0;
        pixel_data[11][70] = 0;
        pixel_data[11][71] = 0;
        pixel_data[11][72] = 0;
        pixel_data[11][73] = 0;
        pixel_data[11][74] = 0;
        pixel_data[11][75] = 0;
        pixel_data[11][76] = 0;
        pixel_data[11][77] = 0;
        pixel_data[11][78] = 0;
        pixel_data[11][79] = 0;
        pixel_data[11][80] = 0;
        pixel_data[11][81] = 0;
        pixel_data[11][82] = 0;
        pixel_data[11][83] = 0;
        pixel_data[11][84] = 0;
        pixel_data[11][85] = 0;
        pixel_data[11][86] = 0;
        pixel_data[11][87] = 0;
        pixel_data[11][88] = 0;
        pixel_data[11][89] = 0;
        pixel_data[11][90] = 0;
        pixel_data[11][91] = 0;
        pixel_data[11][92] = 0;
        pixel_data[11][93] = 0;
        pixel_data[11][94] = 0;
        pixel_data[11][95] = 0;
        pixel_data[11][96] = 0;
        pixel_data[11][97] = 0;
        pixel_data[11][98] = 0;
        pixel_data[11][99] = 0; // y=11
        pixel_data[12][0] = 0;
        pixel_data[12][1] = 0;
        pixel_data[12][2] = 0;
        pixel_data[12][3] = 0;
        pixel_data[12][4] = 0;
        pixel_data[12][5] = 0;
        pixel_data[12][6] = 0;
        pixel_data[12][7] = 0;
        pixel_data[12][8] = 0;
        pixel_data[12][9] = 0;
        pixel_data[12][10] = 0;
        pixel_data[12][11] = 0;
        pixel_data[12][12] = 0;
        pixel_data[12][13] = 0;
        pixel_data[12][14] = 0;
        pixel_data[12][15] = 0;
        pixel_data[12][16] = 0;
        pixel_data[12][17] = 0;
        pixel_data[12][18] = 0;
        pixel_data[12][19] = 0;
        pixel_data[12][20] = 0;
        pixel_data[12][21] = 0;
        pixel_data[12][22] = 0;
        pixel_data[12][23] = 0;
        pixel_data[12][24] = 0;
        pixel_data[12][25] = 0;
        pixel_data[12][26] = 0;
        pixel_data[12][27] = 0;
        pixel_data[12][28] = 0;
        pixel_data[12][29] = 0;
        pixel_data[12][30] = 0;
        pixel_data[12][31] = 0;
        pixel_data[12][32] = 0;
        pixel_data[12][33] = 0;
        pixel_data[12][34] = 0;
        pixel_data[12][35] = 0;
        pixel_data[12][36] = 0;
        pixel_data[12][37] = 0;
        pixel_data[12][38] = 0;
        pixel_data[12][39] = 0;
        pixel_data[12][40] = 0;
        pixel_data[12][41] = 0;
        pixel_data[12][42] = 0;
        pixel_data[12][43] = 0;
        pixel_data[12][44] = 0;
        pixel_data[12][45] = 0;
        pixel_data[12][46] = 0;
        pixel_data[12][47] = 0;
        pixel_data[12][48] = 0;
        pixel_data[12][49] = 0;
        pixel_data[12][50] = 0;
        pixel_data[12][51] = 0;
        pixel_data[12][52] = 0;
        pixel_data[12][53] = 0;
        pixel_data[12][54] = 0;
        pixel_data[12][55] = 0;
        pixel_data[12][56] = 0;
        pixel_data[12][57] = 0;
        pixel_data[12][58] = 0;
        pixel_data[12][59] = 0;
        pixel_data[12][60] = 0;
        pixel_data[12][61] = 0;
        pixel_data[12][62] = 0;
        pixel_data[12][63] = 0;
        pixel_data[12][64] = 0;
        pixel_data[12][65] = 0;
        pixel_data[12][66] = 0;
        pixel_data[12][67] = 0;
        pixel_data[12][68] = 0;
        pixel_data[12][69] = 0;
        pixel_data[12][70] = 0;
        pixel_data[12][71] = 0;
        pixel_data[12][72] = 0;
        pixel_data[12][73] = 0;
        pixel_data[12][74] = 0;
        pixel_data[12][75] = 0;
        pixel_data[12][76] = 0;
        pixel_data[12][77] = 0;
        pixel_data[12][78] = 0;
        pixel_data[12][79] = 0;
        pixel_data[12][80] = 0;
        pixel_data[12][81] = 0;
        pixel_data[12][82] = 0;
        pixel_data[12][83] = 0;
        pixel_data[12][84] = 0;
        pixel_data[12][85] = 0;
        pixel_data[12][86] = 0;
        pixel_data[12][87] = 0;
        pixel_data[12][88] = 0;
        pixel_data[12][89] = 0;
        pixel_data[12][90] = 0;
        pixel_data[12][91] = 0;
        pixel_data[12][92] = 0;
        pixel_data[12][93] = 0;
        pixel_data[12][94] = 0;
        pixel_data[12][95] = 0;
        pixel_data[12][96] = 0;
        pixel_data[12][97] = 0;
        pixel_data[12][98] = 0;
        pixel_data[12][99] = 0; // y=12
        pixel_data[13][0] = 0;
        pixel_data[13][1] = 0;
        pixel_data[13][2] = 0;
        pixel_data[13][3] = 0;
        pixel_data[13][4] = 0;
        pixel_data[13][5] = 0;
        pixel_data[13][6] = 0;
        pixel_data[13][7] = 0;
        pixel_data[13][8] = 0;
        pixel_data[13][9] = 0;
        pixel_data[13][10] = 0;
        pixel_data[13][11] = 0;
        pixel_data[13][12] = 0;
        pixel_data[13][13] = 0;
        pixel_data[13][14] = 0;
        pixel_data[13][15] = 0;
        pixel_data[13][16] = 0;
        pixel_data[13][17] = 0;
        pixel_data[13][18] = 0;
        pixel_data[13][19] = 0;
        pixel_data[13][20] = 0;
        pixel_data[13][21] = 0;
        pixel_data[13][22] = 0;
        pixel_data[13][23] = 0;
        pixel_data[13][24] = 0;
        pixel_data[13][25] = 0;
        pixel_data[13][26] = 0;
        pixel_data[13][27] = 0;
        pixel_data[13][28] = 0;
        pixel_data[13][29] = 0;
        pixel_data[13][30] = 0;
        pixel_data[13][31] = 0;
        pixel_data[13][32] = 0;
        pixel_data[13][33] = 0;
        pixel_data[13][34] = 0;
        pixel_data[13][35] = 0;
        pixel_data[13][36] = 0;
        pixel_data[13][37] = 0;
        pixel_data[13][38] = 0;
        pixel_data[13][39] = 0;
        pixel_data[13][40] = 0;
        pixel_data[13][41] = 0;
        pixel_data[13][42] = 0;
        pixel_data[13][43] = 0;
        pixel_data[13][44] = 0;
        pixel_data[13][45] = 0;
        pixel_data[13][46] = 0;
        pixel_data[13][47] = 0;
        pixel_data[13][48] = 0;
        pixel_data[13][49] = 0;
        pixel_data[13][50] = 0;
        pixel_data[13][51] = 0;
        pixel_data[13][52] = 0;
        pixel_data[13][53] = 0;
        pixel_data[13][54] = 0;
        pixel_data[13][55] = 0;
        pixel_data[13][56] = 0;
        pixel_data[13][57] = 0;
        pixel_data[13][58] = 0;
        pixel_data[13][59] = 0;
        pixel_data[13][60] = 0;
        pixel_data[13][61] = 0;
        pixel_data[13][62] = 0;
        pixel_data[13][63] = 0;
        pixel_data[13][64] = 0;
        pixel_data[13][65] = 0;
        pixel_data[13][66] = 0;
        pixel_data[13][67] = 0;
        pixel_data[13][68] = 0;
        pixel_data[13][69] = 0;
        pixel_data[13][70] = 0;
        pixel_data[13][71] = 0;
        pixel_data[13][72] = 0;
        pixel_data[13][73] = 0;
        pixel_data[13][74] = 0;
        pixel_data[13][75] = 0;
        pixel_data[13][76] = 0;
        pixel_data[13][77] = 0;
        pixel_data[13][78] = 0;
        pixel_data[13][79] = 0;
        pixel_data[13][80] = 0;
        pixel_data[13][81] = 0;
        pixel_data[13][82] = 0;
        pixel_data[13][83] = 0;
        pixel_data[13][84] = 0;
        pixel_data[13][85] = 0;
        pixel_data[13][86] = 0;
        pixel_data[13][87] = 0;
        pixel_data[13][88] = 0;
        pixel_data[13][89] = 0;
        pixel_data[13][90] = 0;
        pixel_data[13][91] = 0;
        pixel_data[13][92] = 0;
        pixel_data[13][93] = 0;
        pixel_data[13][94] = 0;
        pixel_data[13][95] = 0;
        pixel_data[13][96] = 0;
        pixel_data[13][97] = 0;
        pixel_data[13][98] = 0;
        pixel_data[13][99] = 0; // y=13
        pixel_data[14][0] = 0;
        pixel_data[14][1] = 0;
        pixel_data[14][2] = 0;
        pixel_data[14][3] = 0;
        pixel_data[14][4] = 0;
        pixel_data[14][5] = 0;
        pixel_data[14][6] = 0;
        pixel_data[14][7] = 0;
        pixel_data[14][8] = 0;
        pixel_data[14][9] = 0;
        pixel_data[14][10] = 0;
        pixel_data[14][11] = 0;
        pixel_data[14][12] = 0;
        pixel_data[14][13] = 0;
        pixel_data[14][14] = 0;
        pixel_data[14][15] = 0;
        pixel_data[14][16] = 0;
        pixel_data[14][17] = 0;
        pixel_data[14][18] = 0;
        pixel_data[14][19] = 0;
        pixel_data[14][20] = 0;
        pixel_data[14][21] = 0;
        pixel_data[14][22] = 0;
        pixel_data[14][23] = 0;
        pixel_data[14][24] = 0;
        pixel_data[14][25] = 0;
        pixel_data[14][26] = 0;
        pixel_data[14][27] = 0;
        pixel_data[14][28] = 0;
        pixel_data[14][29] = 0;
        pixel_data[14][30] = 0;
        pixel_data[14][31] = 0;
        pixel_data[14][32] = 0;
        pixel_data[14][33] = 0;
        pixel_data[14][34] = 0;
        pixel_data[14][35] = 0;
        pixel_data[14][36] = 0;
        pixel_data[14][37] = 0;
        pixel_data[14][38] = 0;
        pixel_data[14][39] = 0;
        pixel_data[14][40] = 0;
        pixel_data[14][41] = 0;
        pixel_data[14][42] = 0;
        pixel_data[14][43] = 0;
        pixel_data[14][44] = 0;
        pixel_data[14][45] = 0;
        pixel_data[14][46] = 0;
        pixel_data[14][47] = 0;
        pixel_data[14][48] = 0;
        pixel_data[14][49] = 0;
        pixel_data[14][50] = 0;
        pixel_data[14][51] = 0;
        pixel_data[14][52] = 0;
        pixel_data[14][53] = 0;
        pixel_data[14][54] = 0;
        pixel_data[14][55] = 0;
        pixel_data[14][56] = 0;
        pixel_data[14][57] = 0;
        pixel_data[14][58] = 0;
        pixel_data[14][59] = 0;
        pixel_data[14][60] = 0;
        pixel_data[14][61] = 0;
        pixel_data[14][62] = 0;
        pixel_data[14][63] = 0;
        pixel_data[14][64] = 0;
        pixel_data[14][65] = 0;
        pixel_data[14][66] = 0;
        pixel_data[14][67] = 0;
        pixel_data[14][68] = 0;
        pixel_data[14][69] = 0;
        pixel_data[14][70] = 0;
        pixel_data[14][71] = 0;
        pixel_data[14][72] = 0;
        pixel_data[14][73] = 0;
        pixel_data[14][74] = 0;
        pixel_data[14][75] = 0;
        pixel_data[14][76] = 0;
        pixel_data[14][77] = 0;
        pixel_data[14][78] = 0;
        pixel_data[14][79] = 0;
        pixel_data[14][80] = 0;
        pixel_data[14][81] = 0;
        pixel_data[14][82] = 0;
        pixel_data[14][83] = 0;
        pixel_data[14][84] = 0;
        pixel_data[14][85] = 0;
        pixel_data[14][86] = 0;
        pixel_data[14][87] = 0;
        pixel_data[14][88] = 0;
        pixel_data[14][89] = 0;
        pixel_data[14][90] = 0;
        pixel_data[14][91] = 0;
        pixel_data[14][92] = 0;
        pixel_data[14][93] = 0;
        pixel_data[14][94] = 0;
        pixel_data[14][95] = 0;
        pixel_data[14][96] = 0;
        pixel_data[14][97] = 0;
        pixel_data[14][98] = 0;
        pixel_data[14][99] = 0; // y=14
        pixel_data[15][0] = 0;
        pixel_data[15][1] = 0;
        pixel_data[15][2] = 0;
        pixel_data[15][3] = 0;
        pixel_data[15][4] = 0;
        pixel_data[15][5] = 0;
        pixel_data[15][6] = 0;
        pixel_data[15][7] = 0;
        pixel_data[15][8] = 0;
        pixel_data[15][9] = 0;
        pixel_data[15][10] = 0;
        pixel_data[15][11] = 0;
        pixel_data[15][12] = 0;
        pixel_data[15][13] = 0;
        pixel_data[15][14] = 0;
        pixel_data[15][15] = 0;
        pixel_data[15][16] = 0;
        pixel_data[15][17] = 0;
        pixel_data[15][18] = 0;
        pixel_data[15][19] = 0;
        pixel_data[15][20] = 0;
        pixel_data[15][21] = 0;
        pixel_data[15][22] = 0;
        pixel_data[15][23] = 0;
        pixel_data[15][24] = 0;
        pixel_data[15][25] = 0;
        pixel_data[15][26] = 0;
        pixel_data[15][27] = 0;
        pixel_data[15][28] = 0;
        pixel_data[15][29] = 0;
        pixel_data[15][30] = 0;
        pixel_data[15][31] = 0;
        pixel_data[15][32] = 0;
        pixel_data[15][33] = 0;
        pixel_data[15][34] = 0;
        pixel_data[15][35] = 0;
        pixel_data[15][36] = 0;
        pixel_data[15][37] = 0;
        pixel_data[15][38] = 0;
        pixel_data[15][39] = 0;
        pixel_data[15][40] = 0;
        pixel_data[15][41] = 0;
        pixel_data[15][42] = 0;
        pixel_data[15][43] = 0;
        pixel_data[15][44] = 0;
        pixel_data[15][45] = 0;
        pixel_data[15][46] = 0;
        pixel_data[15][47] = 0;
        pixel_data[15][48] = 0;
        pixel_data[15][49] = 0;
        pixel_data[15][50] = 0;
        pixel_data[15][51] = 0;
        pixel_data[15][52] = 0;
        pixel_data[15][53] = 0;
        pixel_data[15][54] = 0;
        pixel_data[15][55] = 0;
        pixel_data[15][56] = 0;
        pixel_data[15][57] = 0;
        pixel_data[15][58] = 0;
        pixel_data[15][59] = 0;
        pixel_data[15][60] = 0;
        pixel_data[15][61] = 0;
        pixel_data[15][62] = 0;
        pixel_data[15][63] = 0;
        pixel_data[15][64] = 0;
        pixel_data[15][65] = 0;
        pixel_data[15][66] = 0;
        pixel_data[15][67] = 0;
        pixel_data[15][68] = 0;
        pixel_data[15][69] = 0;
        pixel_data[15][70] = 0;
        pixel_data[15][71] = 0;
        pixel_data[15][72] = 0;
        pixel_data[15][73] = 0;
        pixel_data[15][74] = 0;
        pixel_data[15][75] = 0;
        pixel_data[15][76] = 0;
        pixel_data[15][77] = 0;
        pixel_data[15][78] = 0;
        pixel_data[15][79] = 0;
        pixel_data[15][80] = 0;
        pixel_data[15][81] = 0;
        pixel_data[15][82] = 0;
        pixel_data[15][83] = 0;
        pixel_data[15][84] = 0;
        pixel_data[15][85] = 0;
        pixel_data[15][86] = 0;
        pixel_data[15][87] = 0;
        pixel_data[15][88] = 0;
        pixel_data[15][89] = 0;
        pixel_data[15][90] = 0;
        pixel_data[15][91] = 0;
        pixel_data[15][92] = 0;
        pixel_data[15][93] = 0;
        pixel_data[15][94] = 0;
        pixel_data[15][95] = 0;
        pixel_data[15][96] = 0;
        pixel_data[15][97] = 0;
        pixel_data[15][98] = 0;
        pixel_data[15][99] = 0; // y=15
        pixel_data[16][0] = 0;
        pixel_data[16][1] = 0;
        pixel_data[16][2] = 0;
        pixel_data[16][3] = 0;
        pixel_data[16][4] = 0;
        pixel_data[16][5] = 0;
        pixel_data[16][6] = 0;
        pixel_data[16][7] = 0;
        pixel_data[16][8] = 0;
        pixel_data[16][9] = 0;
        pixel_data[16][10] = 0;
        pixel_data[16][11] = 0;
        pixel_data[16][12] = 0;
        pixel_data[16][13] = 0;
        pixel_data[16][14] = 0;
        pixel_data[16][15] = 0;
        pixel_data[16][16] = 0;
        pixel_data[16][17] = 0;
        pixel_data[16][18] = 0;
        pixel_data[16][19] = 0;
        pixel_data[16][20] = 0;
        pixel_data[16][21] = 0;
        pixel_data[16][22] = 0;
        pixel_data[16][23] = 0;
        pixel_data[16][24] = 0;
        pixel_data[16][25] = 0;
        pixel_data[16][26] = 0;
        pixel_data[16][27] = 0;
        pixel_data[16][28] = 0;
        pixel_data[16][29] = 0;
        pixel_data[16][30] = 0;
        pixel_data[16][31] = 0;
        pixel_data[16][32] = 0;
        pixel_data[16][33] = 0;
        pixel_data[16][34] = 0;
        pixel_data[16][35] = 0;
        pixel_data[16][36] = 0;
        pixel_data[16][37] = 0;
        pixel_data[16][38] = 0;
        pixel_data[16][39] = 0;
        pixel_data[16][40] = 0;
        pixel_data[16][41] = 0;
        pixel_data[16][42] = 0;
        pixel_data[16][43] = 0;
        pixel_data[16][44] = 0;
        pixel_data[16][45] = 0;
        pixel_data[16][46] = 0;
        pixel_data[16][47] = 0;
        pixel_data[16][48] = 0;
        pixel_data[16][49] = 0;
        pixel_data[16][50] = 0;
        pixel_data[16][51] = 0;
        pixel_data[16][52] = 0;
        pixel_data[16][53] = 0;
        pixel_data[16][54] = 0;
        pixel_data[16][55] = 0;
        pixel_data[16][56] = 0;
        pixel_data[16][57] = 0;
        pixel_data[16][58] = 0;
        pixel_data[16][59] = 0;
        pixel_data[16][60] = 0;
        pixel_data[16][61] = 0;
        pixel_data[16][62] = 0;
        pixel_data[16][63] = 0;
        pixel_data[16][64] = 0;
        pixel_data[16][65] = 0;
        pixel_data[16][66] = 0;
        pixel_data[16][67] = 0;
        pixel_data[16][68] = 0;
        pixel_data[16][69] = 0;
        pixel_data[16][70] = 0;
        pixel_data[16][71] = 0;
        pixel_data[16][72] = 0;
        pixel_data[16][73] = 0;
        pixel_data[16][74] = 0;
        pixel_data[16][75] = 0;
        pixel_data[16][76] = 0;
        pixel_data[16][77] = 0;
        pixel_data[16][78] = 0;
        pixel_data[16][79] = 0;
        pixel_data[16][80] = 0;
        pixel_data[16][81] = 0;
        pixel_data[16][82] = 0;
        pixel_data[16][83] = 0;
        pixel_data[16][84] = 0;
        pixel_data[16][85] = 0;
        pixel_data[16][86] = 0;
        pixel_data[16][87] = 0;
        pixel_data[16][88] = 0;
        pixel_data[16][89] = 0;
        pixel_data[16][90] = 0;
        pixel_data[16][91] = 0;
        pixel_data[16][92] = 0;
        pixel_data[16][93] = 0;
        pixel_data[16][94] = 0;
        pixel_data[16][95] = 0;
        pixel_data[16][96] = 0;
        pixel_data[16][97] = 0;
        pixel_data[16][98] = 0;
        pixel_data[16][99] = 0; // y=16
        pixel_data[17][0] = 0;
        pixel_data[17][1] = 0;
        pixel_data[17][2] = 0;
        pixel_data[17][3] = 0;
        pixel_data[17][4] = 0;
        pixel_data[17][5] = 0;
        pixel_data[17][6] = 0;
        pixel_data[17][7] = 0;
        pixel_data[17][8] = 0;
        pixel_data[17][9] = 0;
        pixel_data[17][10] = 0;
        pixel_data[17][11] = 0;
        pixel_data[17][12] = 0;
        pixel_data[17][13] = 0;
        pixel_data[17][14] = 0;
        pixel_data[17][15] = 0;
        pixel_data[17][16] = 0;
        pixel_data[17][17] = 0;
        pixel_data[17][18] = 0;
        pixel_data[17][19] = 0;
        pixel_data[17][20] = 0;
        pixel_data[17][21] = 0;
        pixel_data[17][22] = 0;
        pixel_data[17][23] = 0;
        pixel_data[17][24] = 0;
        pixel_data[17][25] = 0;
        pixel_data[17][26] = 0;
        pixel_data[17][27] = 0;
        pixel_data[17][28] = 0;
        pixel_data[17][29] = 0;
        pixel_data[17][30] = 0;
        pixel_data[17][31] = 0;
        pixel_data[17][32] = 0;
        pixel_data[17][33] = 0;
        pixel_data[17][34] = 0;
        pixel_data[17][35] = 0;
        pixel_data[17][36] = 0;
        pixel_data[17][37] = 0;
        pixel_data[17][38] = 0;
        pixel_data[17][39] = 0;
        pixel_data[17][40] = 0;
        pixel_data[17][41] = 0;
        pixel_data[17][42] = 0;
        pixel_data[17][43] = 0;
        pixel_data[17][44] = 0;
        pixel_data[17][45] = 0;
        pixel_data[17][46] = 0;
        pixel_data[17][47] = 0;
        pixel_data[17][48] = 0;
        pixel_data[17][49] = 0;
        pixel_data[17][50] = 0;
        pixel_data[17][51] = 0;
        pixel_data[17][52] = 0;
        pixel_data[17][53] = 0;
        pixel_data[17][54] = 0;
        pixel_data[17][55] = 0;
        pixel_data[17][56] = 0;
        pixel_data[17][57] = 0;
        pixel_data[17][58] = 0;
        pixel_data[17][59] = 0;
        pixel_data[17][60] = 0;
        pixel_data[17][61] = 0;
        pixel_data[17][62] = 0;
        pixel_data[17][63] = 0;
        pixel_data[17][64] = 0;
        pixel_data[17][65] = 0;
        pixel_data[17][66] = 0;
        pixel_data[17][67] = 0;
        pixel_data[17][68] = 0;
        pixel_data[17][69] = 0;
        pixel_data[17][70] = 0;
        pixel_data[17][71] = 0;
        pixel_data[17][72] = 0;
        pixel_data[17][73] = 0;
        pixel_data[17][74] = 0;
        pixel_data[17][75] = 0;
        pixel_data[17][76] = 0;
        pixel_data[17][77] = 0;
        pixel_data[17][78] = 0;
        pixel_data[17][79] = 0;
        pixel_data[17][80] = 0;
        pixel_data[17][81] = 0;
        pixel_data[17][82] = 0;
        pixel_data[17][83] = 0;
        pixel_data[17][84] = 0;
        pixel_data[17][85] = 0;
        pixel_data[17][86] = 0;
        pixel_data[17][87] = 0;
        pixel_data[17][88] = 0;
        pixel_data[17][89] = 0;
        pixel_data[17][90] = 0;
        pixel_data[17][91] = 0;
        pixel_data[17][92] = 0;
        pixel_data[17][93] = 0;
        pixel_data[17][94] = 0;
        pixel_data[17][95] = 0;
        pixel_data[17][96] = 0;
        pixel_data[17][97] = 0;
        pixel_data[17][98] = 0;
        pixel_data[17][99] = 0; // y=17
        pixel_data[18][0] = 0;
        pixel_data[18][1] = 0;
        pixel_data[18][2] = 0;
        pixel_data[18][3] = 0;
        pixel_data[18][4] = 0;
        pixel_data[18][5] = 0;
        pixel_data[18][6] = 0;
        pixel_data[18][7] = 0;
        pixel_data[18][8] = 0;
        pixel_data[18][9] = 0;
        pixel_data[18][10] = 0;
        pixel_data[18][11] = 0;
        pixel_data[18][12] = 0;
        pixel_data[18][13] = 0;
        pixel_data[18][14] = 0;
        pixel_data[18][15] = 0;
        pixel_data[18][16] = 0;
        pixel_data[18][17] = 0;
        pixel_data[18][18] = 0;
        pixel_data[18][19] = 0;
        pixel_data[18][20] = 0;
        pixel_data[18][21] = 0;
        pixel_data[18][22] = 0;
        pixel_data[18][23] = 0;
        pixel_data[18][24] = 0;
        pixel_data[18][25] = 0;
        pixel_data[18][26] = 0;
        pixel_data[18][27] = 0;
        pixel_data[18][28] = 0;
        pixel_data[18][29] = 0;
        pixel_data[18][30] = 0;
        pixel_data[18][31] = 0;
        pixel_data[18][32] = 0;
        pixel_data[18][33] = 0;
        pixel_data[18][34] = 0;
        pixel_data[18][35] = 0;
        pixel_data[18][36] = 0;
        pixel_data[18][37] = 0;
        pixel_data[18][38] = 0;
        pixel_data[18][39] = 0;
        pixel_data[18][40] = 0;
        pixel_data[18][41] = 0;
        pixel_data[18][42] = 0;
        pixel_data[18][43] = 0;
        pixel_data[18][44] = 0;
        pixel_data[18][45] = 0;
        pixel_data[18][46] = 0;
        pixel_data[18][47] = 0;
        pixel_data[18][48] = 0;
        pixel_data[18][49] = 0;
        pixel_data[18][50] = 0;
        pixel_data[18][51] = 0;
        pixel_data[18][52] = 0;
        pixel_data[18][53] = 0;
        pixel_data[18][54] = 0;
        pixel_data[18][55] = 0;
        pixel_data[18][56] = 0;
        pixel_data[18][57] = 0;
        pixel_data[18][58] = 0;
        pixel_data[18][59] = 0;
        pixel_data[18][60] = 0;
        pixel_data[18][61] = 0;
        pixel_data[18][62] = 0;
        pixel_data[18][63] = 0;
        pixel_data[18][64] = 0;
        pixel_data[18][65] = 0;
        pixel_data[18][66] = 0;
        pixel_data[18][67] = 0;
        pixel_data[18][68] = 0;
        pixel_data[18][69] = 0;
        pixel_data[18][70] = 0;
        pixel_data[18][71] = 0;
        pixel_data[18][72] = 0;
        pixel_data[18][73] = 0;
        pixel_data[18][74] = 0;
        pixel_data[18][75] = 0;
        pixel_data[18][76] = 0;
        pixel_data[18][77] = 0;
        pixel_data[18][78] = 0;
        pixel_data[18][79] = 0;
        pixel_data[18][80] = 0;
        pixel_data[18][81] = 0;
        pixel_data[18][82] = 0;
        pixel_data[18][83] = 0;
        pixel_data[18][84] = 0;
        pixel_data[18][85] = 0;
        pixel_data[18][86] = 0;
        pixel_data[18][87] = 0;
        pixel_data[18][88] = 0;
        pixel_data[18][89] = 0;
        pixel_data[18][90] = 0;
        pixel_data[18][91] = 0;
        pixel_data[18][92] = 0;
        pixel_data[18][93] = 0;
        pixel_data[18][94] = 0;
        pixel_data[18][95] = 0;
        pixel_data[18][96] = 0;
        pixel_data[18][97] = 0;
        pixel_data[18][98] = 0;
        pixel_data[18][99] = 0; // y=18
        pixel_data[19][0] = 0;
        pixel_data[19][1] = 0;
        pixel_data[19][2] = 0;
        pixel_data[19][3] = 0;
        pixel_data[19][4] = 0;
        pixel_data[19][5] = 0;
        pixel_data[19][6] = 0;
        pixel_data[19][7] = 0;
        pixel_data[19][8] = 0;
        pixel_data[19][9] = 0;
        pixel_data[19][10] = 0;
        pixel_data[19][11] = 0;
        pixel_data[19][12] = 0;
        pixel_data[19][13] = 0;
        pixel_data[19][14] = 0;
        pixel_data[19][15] = 0;
        pixel_data[19][16] = 0;
        pixel_data[19][17] = 0;
        pixel_data[19][18] = 0;
        pixel_data[19][19] = 0;
        pixel_data[19][20] = 0;
        pixel_data[19][21] = 0;
        pixel_data[19][22] = 0;
        pixel_data[19][23] = 0;
        pixel_data[19][24] = 0;
        pixel_data[19][25] = 0;
        pixel_data[19][26] = 0;
        pixel_data[19][27] = 0;
        pixel_data[19][28] = 0;
        pixel_data[19][29] = 0;
        pixel_data[19][30] = 0;
        pixel_data[19][31] = 0;
        pixel_data[19][32] = 0;
        pixel_data[19][33] = 0;
        pixel_data[19][34] = 0;
        pixel_data[19][35] = 0;
        pixel_data[19][36] = 0;
        pixel_data[19][37] = 0;
        pixel_data[19][38] = 0;
        pixel_data[19][39] = 0;
        pixel_data[19][40] = 0;
        pixel_data[19][41] = 0;
        pixel_data[19][42] = 0;
        pixel_data[19][43] = 0;
        pixel_data[19][44] = 0;
        pixel_data[19][45] = 0;
        pixel_data[19][46] = 0;
        pixel_data[19][47] = 0;
        pixel_data[19][48] = 0;
        pixel_data[19][49] = 0;
        pixel_data[19][50] = 0;
        pixel_data[19][51] = 0;
        pixel_data[19][52] = 0;
        pixel_data[19][53] = 0;
        pixel_data[19][54] = 0;
        pixel_data[19][55] = 0;
        pixel_data[19][56] = 0;
        pixel_data[19][57] = 0;
        pixel_data[19][58] = 0;
        pixel_data[19][59] = 0;
        pixel_data[19][60] = 0;
        pixel_data[19][61] = 0;
        pixel_data[19][62] = 0;
        pixel_data[19][63] = 0;
        pixel_data[19][64] = 0;
        pixel_data[19][65] = 0;
        pixel_data[19][66] = 0;
        pixel_data[19][67] = 0;
        pixel_data[19][68] = 0;
        pixel_data[19][69] = 0;
        pixel_data[19][70] = 0;
        pixel_data[19][71] = 0;
        pixel_data[19][72] = 0;
        pixel_data[19][73] = 0;
        pixel_data[19][74] = 0;
        pixel_data[19][75] = 0;
        pixel_data[19][76] = 0;
        pixel_data[19][77] = 0;
        pixel_data[19][78] = 0;
        pixel_data[19][79] = 0;
        pixel_data[19][80] = 0;
        pixel_data[19][81] = 0;
        pixel_data[19][82] = 0;
        pixel_data[19][83] = 0;
        pixel_data[19][84] = 0;
        pixel_data[19][85] = 0;
        pixel_data[19][86] = 0;
        pixel_data[19][87] = 0;
        pixel_data[19][88] = 0;
        pixel_data[19][89] = 0;
        pixel_data[19][90] = 0;
        pixel_data[19][91] = 0;
        pixel_data[19][92] = 0;
        pixel_data[19][93] = 0;
        pixel_data[19][94] = 0;
        pixel_data[19][95] = 0;
        pixel_data[19][96] = 0;
        pixel_data[19][97] = 0;
        pixel_data[19][98] = 0;
        pixel_data[19][99] = 0; // y=19
        pixel_data[20][0] = 0;
        pixel_data[20][1] = 0;
        pixel_data[20][2] = 0;
        pixel_data[20][3] = 0;
        pixel_data[20][4] = 0;
        pixel_data[20][5] = 0;
        pixel_data[20][6] = 0;
        pixel_data[20][7] = 0;
        pixel_data[20][8] = 0;
        pixel_data[20][9] = 0;
        pixel_data[20][10] = 0;
        pixel_data[20][11] = 0;
        pixel_data[20][12] = 0;
        pixel_data[20][13] = 0;
        pixel_data[20][14] = 0;
        pixel_data[20][15] = 0;
        pixel_data[20][16] = 0;
        pixel_data[20][17] = 0;
        pixel_data[20][18] = 0;
        pixel_data[20][19] = 0;
        pixel_data[20][20] = 0;
        pixel_data[20][21] = 0;
        pixel_data[20][22] = 0;
        pixel_data[20][23] = 0;
        pixel_data[20][24] = 0;
        pixel_data[20][25] = 0;
        pixel_data[20][26] = 0;
        pixel_data[20][27] = 0;
        pixel_data[20][28] = 0;
        pixel_data[20][29] = 0;
        pixel_data[20][30] = 0;
        pixel_data[20][31] = 0;
        pixel_data[20][32] = 0;
        pixel_data[20][33] = 0;
        pixel_data[20][34] = 0;
        pixel_data[20][35] = 0;
        pixel_data[20][36] = 0;
        pixel_data[20][37] = 0;
        pixel_data[20][38] = 0;
        pixel_data[20][39] = 0;
        pixel_data[20][40] = 0;
        pixel_data[20][41] = 0;
        pixel_data[20][42] = 0;
        pixel_data[20][43] = 0;
        pixel_data[20][44] = 0;
        pixel_data[20][45] = 0;
        pixel_data[20][46] = 0;
        pixel_data[20][47] = 0;
        pixel_data[20][48] = 0;
        pixel_data[20][49] = 0;
        pixel_data[20][50] = 0;
        pixel_data[20][51] = 0;
        pixel_data[20][52] = 0;
        pixel_data[20][53] = 0;
        pixel_data[20][54] = 0;
        pixel_data[20][55] = 0;
        pixel_data[20][56] = 0;
        pixel_data[20][57] = 0;
        pixel_data[20][58] = 0;
        pixel_data[20][59] = 0;
        pixel_data[20][60] = 0;
        pixel_data[20][61] = 0;
        pixel_data[20][62] = 0;
        pixel_data[20][63] = 0;
        pixel_data[20][64] = 0;
        pixel_data[20][65] = 0;
        pixel_data[20][66] = 0;
        pixel_data[20][67] = 0;
        pixel_data[20][68] = 0;
        pixel_data[20][69] = 0;
        pixel_data[20][70] = 0;
        pixel_data[20][71] = 0;
        pixel_data[20][72] = 0;
        pixel_data[20][73] = 0;
        pixel_data[20][74] = 0;
        pixel_data[20][75] = 0;
        pixel_data[20][76] = 0;
        pixel_data[20][77] = 0;
        pixel_data[20][78] = 0;
        pixel_data[20][79] = 0;
        pixel_data[20][80] = 0;
        pixel_data[20][81] = 0;
        pixel_data[20][82] = 0;
        pixel_data[20][83] = 0;
        pixel_data[20][84] = 0;
        pixel_data[20][85] = 0;
        pixel_data[20][86] = 0;
        pixel_data[20][87] = 0;
        pixel_data[20][88] = 0;
        pixel_data[20][89] = 0;
        pixel_data[20][90] = 0;
        pixel_data[20][91] = 0;
        pixel_data[20][92] = 0;
        pixel_data[20][93] = 0;
        pixel_data[20][94] = 0;
        pixel_data[20][95] = 0;
        pixel_data[20][96] = 0;
        pixel_data[20][97] = 0;
        pixel_data[20][98] = 0;
        pixel_data[20][99] = 0; // y=20
        pixel_data[21][0] = 0;
        pixel_data[21][1] = 0;
        pixel_data[21][2] = 0;
        pixel_data[21][3] = 0;
        pixel_data[21][4] = 0;
        pixel_data[21][5] = 0;
        pixel_data[21][6] = 0;
        pixel_data[21][7] = 0;
        pixel_data[21][8] = 0;
        pixel_data[21][9] = 0;
        pixel_data[21][10] = 0;
        pixel_data[21][11] = 0;
        pixel_data[21][12] = 0;
        pixel_data[21][13] = 0;
        pixel_data[21][14] = 0;
        pixel_data[21][15] = 0;
        pixel_data[21][16] = 0;
        pixel_data[21][17] = 0;
        pixel_data[21][18] = 0;
        pixel_data[21][19] = 0;
        pixel_data[21][20] = 0;
        pixel_data[21][21] = 0;
        pixel_data[21][22] = 0;
        pixel_data[21][23] = 0;
        pixel_data[21][24] = 0;
        pixel_data[21][25] = 0;
        pixel_data[21][26] = 0;
        pixel_data[21][27] = 0;
        pixel_data[21][28] = 0;
        pixel_data[21][29] = 0;
        pixel_data[21][30] = 0;
        pixel_data[21][31] = 0;
        pixel_data[21][32] = 0;
        pixel_data[21][33] = 0;
        pixel_data[21][34] = 0;
        pixel_data[21][35] = 0;
        pixel_data[21][36] = 0;
        pixel_data[21][37] = 0;
        pixel_data[21][38] = 0;
        pixel_data[21][39] = 0;
        pixel_data[21][40] = 0;
        pixel_data[21][41] = 0;
        pixel_data[21][42] = 0;
        pixel_data[21][43] = 0;
        pixel_data[21][44] = 0;
        pixel_data[21][45] = 0;
        pixel_data[21][46] = 0;
        pixel_data[21][47] = 0;
        pixel_data[21][48] = 0;
        pixel_data[21][49] = 0;
        pixel_data[21][50] = 0;
        pixel_data[21][51] = 0;
        pixel_data[21][52] = 0;
        pixel_data[21][53] = 0;
        pixel_data[21][54] = 0;
        pixel_data[21][55] = 0;
        pixel_data[21][56] = 0;
        pixel_data[21][57] = 0;
        pixel_data[21][58] = 0;
        pixel_data[21][59] = 0;
        pixel_data[21][60] = 0;
        pixel_data[21][61] = 0;
        pixel_data[21][62] = 0;
        pixel_data[21][63] = 0;
        pixel_data[21][64] = 0;
        pixel_data[21][65] = 0;
        pixel_data[21][66] = 0;
        pixel_data[21][67] = 0;
        pixel_data[21][68] = 0;
        pixel_data[21][69] = 0;
        pixel_data[21][70] = 0;
        pixel_data[21][71] = 0;
        pixel_data[21][72] = 0;
        pixel_data[21][73] = 0;
        pixel_data[21][74] = 0;
        pixel_data[21][75] = 0;
        pixel_data[21][76] = 0;
        pixel_data[21][77] = 0;
        pixel_data[21][78] = 0;
        pixel_data[21][79] = 0;
        pixel_data[21][80] = 0;
        pixel_data[21][81] = 0;
        pixel_data[21][82] = 0;
        pixel_data[21][83] = 0;
        pixel_data[21][84] = 0;
        pixel_data[21][85] = 0;
        pixel_data[21][86] = 0;
        pixel_data[21][87] = 0;
        pixel_data[21][88] = 0;
        pixel_data[21][89] = 0;
        pixel_data[21][90] = 0;
        pixel_data[21][91] = 0;
        pixel_data[21][92] = 0;
        pixel_data[21][93] = 0;
        pixel_data[21][94] = 0;
        pixel_data[21][95] = 0;
        pixel_data[21][96] = 0;
        pixel_data[21][97] = 0;
        pixel_data[21][98] = 0;
        pixel_data[21][99] = 0; // y=21
        pixel_data[22][0] = 0;
        pixel_data[22][1] = 0;
        pixel_data[22][2] = 0;
        pixel_data[22][3] = 0;
        pixel_data[22][4] = 0;
        pixel_data[22][5] = 0;
        pixel_data[22][6] = 0;
        pixel_data[22][7] = 0;
        pixel_data[22][8] = 0;
        pixel_data[22][9] = 0;
        pixel_data[22][10] = 0;
        pixel_data[22][11] = 0;
        pixel_data[22][12] = 0;
        pixel_data[22][13] = 0;
        pixel_data[22][14] = 0;
        pixel_data[22][15] = 0;
        pixel_data[22][16] = 0;
        pixel_data[22][17] = 0;
        pixel_data[22][18] = 0;
        pixel_data[22][19] = 0;
        pixel_data[22][20] = 0;
        pixel_data[22][21] = 0;
        pixel_data[22][22] = 0;
        pixel_data[22][23] = 0;
        pixel_data[22][24] = 0;
        pixel_data[22][25] = 0;
        pixel_data[22][26] = 0;
        pixel_data[22][27] = 0;
        pixel_data[22][28] = 0;
        pixel_data[22][29] = 0;
        pixel_data[22][30] = 0;
        pixel_data[22][31] = 0;
        pixel_data[22][32] = 0;
        pixel_data[22][33] = 0;
        pixel_data[22][34] = 0;
        pixel_data[22][35] = 0;
        pixel_data[22][36] = 0;
        pixel_data[22][37] = 0;
        pixel_data[22][38] = 0;
        pixel_data[22][39] = 0;
        pixel_data[22][40] = 0;
        pixel_data[22][41] = 0;
        pixel_data[22][42] = 0;
        pixel_data[22][43] = 0;
        pixel_data[22][44] = 0;
        pixel_data[22][45] = 0;
        pixel_data[22][46] = 0;
        pixel_data[22][47] = 0;
        pixel_data[22][48] = 0;
        pixel_data[22][49] = 0;
        pixel_data[22][50] = 0;
        pixel_data[22][51] = 0;
        pixel_data[22][52] = 0;
        pixel_data[22][53] = 0;
        pixel_data[22][54] = 0;
        pixel_data[22][55] = 0;
        pixel_data[22][56] = 0;
        pixel_data[22][57] = 0;
        pixel_data[22][58] = 0;
        pixel_data[22][59] = 0;
        pixel_data[22][60] = 0;
        pixel_data[22][61] = 0;
        pixel_data[22][62] = 0;
        pixel_data[22][63] = 0;
        pixel_data[22][64] = 0;
        pixel_data[22][65] = 0;
        pixel_data[22][66] = 0;
        pixel_data[22][67] = 0;
        pixel_data[22][68] = 0;
        pixel_data[22][69] = 0;
        pixel_data[22][70] = 0;
        pixel_data[22][71] = 0;
        pixel_data[22][72] = 0;
        pixel_data[22][73] = 0;
        pixel_data[22][74] = 0;
        pixel_data[22][75] = 0;
        pixel_data[22][76] = 0;
        pixel_data[22][77] = 0;
        pixel_data[22][78] = 0;
        pixel_data[22][79] = 0;
        pixel_data[22][80] = 0;
        pixel_data[22][81] = 0;
        pixel_data[22][82] = 0;
        pixel_data[22][83] = 0;
        pixel_data[22][84] = 0;
        pixel_data[22][85] = 0;
        pixel_data[22][86] = 0;
        pixel_data[22][87] = 0;
        pixel_data[22][88] = 0;
        pixel_data[22][89] = 0;
        pixel_data[22][90] = 0;
        pixel_data[22][91] = 0;
        pixel_data[22][92] = 0;
        pixel_data[22][93] = 0;
        pixel_data[22][94] = 0;
        pixel_data[22][95] = 0;
        pixel_data[22][96] = 0;
        pixel_data[22][97] = 0;
        pixel_data[22][98] = 0;
        pixel_data[22][99] = 0; // y=22
        pixel_data[23][0] = 0;
        pixel_data[23][1] = 0;
        pixel_data[23][2] = 0;
        pixel_data[23][3] = 0;
        pixel_data[23][4] = 0;
        pixel_data[23][5] = 0;
        pixel_data[23][6] = 0;
        pixel_data[23][7] = 0;
        pixel_data[23][8] = 0;
        pixel_data[23][9] = 0;
        pixel_data[23][10] = 0;
        pixel_data[23][11] = 0;
        pixel_data[23][12] = 0;
        pixel_data[23][13] = 0;
        pixel_data[23][14] = 0;
        pixel_data[23][15] = 0;
        pixel_data[23][16] = 0;
        pixel_data[23][17] = 0;
        pixel_data[23][18] = 0;
        pixel_data[23][19] = 0;
        pixel_data[23][20] = 0;
        pixel_data[23][21] = 0;
        pixel_data[23][22] = 0;
        pixel_data[23][23] = 0;
        pixel_data[23][24] = 0;
        pixel_data[23][25] = 0;
        pixel_data[23][26] = 0;
        pixel_data[23][27] = 0;
        pixel_data[23][28] = 0;
        pixel_data[23][29] = 0;
        pixel_data[23][30] = 0;
        pixel_data[23][31] = 0;
        pixel_data[23][32] = 0;
        pixel_data[23][33] = 0;
        pixel_data[23][34] = 0;
        pixel_data[23][35] = 0;
        pixel_data[23][36] = 0;
        pixel_data[23][37] = 0;
        pixel_data[23][38] = 0;
        pixel_data[23][39] = 0;
        pixel_data[23][40] = 0;
        pixel_data[23][41] = 0;
        pixel_data[23][42] = 0;
        pixel_data[23][43] = 0;
        pixel_data[23][44] = 0;
        pixel_data[23][45] = 0;
        pixel_data[23][46] = 0;
        pixel_data[23][47] = 0;
        pixel_data[23][48] = 0;
        pixel_data[23][49] = 0;
        pixel_data[23][50] = 0;
        pixel_data[23][51] = 0;
        pixel_data[23][52] = 0;
        pixel_data[23][53] = 0;
        pixel_data[23][54] = 0;
        pixel_data[23][55] = 0;
        pixel_data[23][56] = 0;
        pixel_data[23][57] = 0;
        pixel_data[23][58] = 0;
        pixel_data[23][59] = 0;
        pixel_data[23][60] = 0;
        pixel_data[23][61] = 0;
        pixel_data[23][62] = 0;
        pixel_data[23][63] = 0;
        pixel_data[23][64] = 0;
        pixel_data[23][65] = 0;
        pixel_data[23][66] = 0;
        pixel_data[23][67] = 0;
        pixel_data[23][68] = 0;
        pixel_data[23][69] = 0;
        pixel_data[23][70] = 0;
        pixel_data[23][71] = 0;
        pixel_data[23][72] = 0;
        pixel_data[23][73] = 0;
        pixel_data[23][74] = 0;
        pixel_data[23][75] = 0;
        pixel_data[23][76] = 0;
        pixel_data[23][77] = 0;
        pixel_data[23][78] = 0;
        pixel_data[23][79] = 0;
        pixel_data[23][80] = 0;
        pixel_data[23][81] = 0;
        pixel_data[23][82] = 0;
        pixel_data[23][83] = 0;
        pixel_data[23][84] = 0;
        pixel_data[23][85] = 0;
        pixel_data[23][86] = 0;
        pixel_data[23][87] = 0;
        pixel_data[23][88] = 0;
        pixel_data[23][89] = 0;
        pixel_data[23][90] = 0;
        pixel_data[23][91] = 0;
        pixel_data[23][92] = 0;
        pixel_data[23][93] = 0;
        pixel_data[23][94] = 0;
        pixel_data[23][95] = 0;
        pixel_data[23][96] = 0;
        pixel_data[23][97] = 0;
        pixel_data[23][98] = 0;
        pixel_data[23][99] = 0; // y=23
        pixel_data[24][0] = 0;
        pixel_data[24][1] = 0;
        pixel_data[24][2] = 0;
        pixel_data[24][3] = 0;
        pixel_data[24][4] = 0;
        pixel_data[24][5] = 0;
        pixel_data[24][6] = 0;
        pixel_data[24][7] = 0;
        pixel_data[24][8] = 0;
        pixel_data[24][9] = 0;
        pixel_data[24][10] = 0;
        pixel_data[24][11] = 0;
        pixel_data[24][12] = 0;
        pixel_data[24][13] = 0;
        pixel_data[24][14] = 0;
        pixel_data[24][15] = 0;
        pixel_data[24][16] = 0;
        pixel_data[24][17] = 0;
        pixel_data[24][18] = 0;
        pixel_data[24][19] = 0;
        pixel_data[24][20] = 0;
        pixel_data[24][21] = 0;
        pixel_data[24][22] = 0;
        pixel_data[24][23] = 0;
        pixel_data[24][24] = 0;
        pixel_data[24][25] = 0;
        pixel_data[24][26] = 0;
        pixel_data[24][27] = 0;
        pixel_data[24][28] = 0;
        pixel_data[24][29] = 0;
        pixel_data[24][30] = 0;
        pixel_data[24][31] = 0;
        pixel_data[24][32] = 0;
        pixel_data[24][33] = 0;
        pixel_data[24][34] = 0;
        pixel_data[24][35] = 0;
        pixel_data[24][36] = 0;
        pixel_data[24][37] = 0;
        pixel_data[24][38] = 0;
        pixel_data[24][39] = 0;
        pixel_data[24][40] = 0;
        pixel_data[24][41] = 0;
        pixel_data[24][42] = 0;
        pixel_data[24][43] = 0;
        pixel_data[24][44] = 0;
        pixel_data[24][45] = 0;
        pixel_data[24][46] = 0;
        pixel_data[24][47] = 0;
        pixel_data[24][48] = 0;
        pixel_data[24][49] = 0;
        pixel_data[24][50] = 0;
        pixel_data[24][51] = 0;
        pixel_data[24][52] = 0;
        pixel_data[24][53] = 0;
        pixel_data[24][54] = 0;
        pixel_data[24][55] = 0;
        pixel_data[24][56] = 0;
        pixel_data[24][57] = 0;
        pixel_data[24][58] = 0;
        pixel_data[24][59] = 0;
        pixel_data[24][60] = 0;
        pixel_data[24][61] = 0;
        pixel_data[24][62] = 0;
        pixel_data[24][63] = 0;
        pixel_data[24][64] = 0;
        pixel_data[24][65] = 0;
        pixel_data[24][66] = 0;
        pixel_data[24][67] = 0;
        pixel_data[24][68] = 0;
        pixel_data[24][69] = 0;
        pixel_data[24][70] = 0;
        pixel_data[24][71] = 0;
        pixel_data[24][72] = 0;
        pixel_data[24][73] = 0;
        pixel_data[24][74] = 0;
        pixel_data[24][75] = 0;
        pixel_data[24][76] = 0;
        pixel_data[24][77] = 0;
        pixel_data[24][78] = 0;
        pixel_data[24][79] = 0;
        pixel_data[24][80] = 0;
        pixel_data[24][81] = 0;
        pixel_data[24][82] = 0;
        pixel_data[24][83] = 0;
        pixel_data[24][84] = 0;
        pixel_data[24][85] = 0;
        pixel_data[24][86] = 0;
        pixel_data[24][87] = 0;
        pixel_data[24][88] = 0;
        pixel_data[24][89] = 0;
        pixel_data[24][90] = 0;
        pixel_data[24][91] = 0;
        pixel_data[24][92] = 0;
        pixel_data[24][93] = 0;
        pixel_data[24][94] = 0;
        pixel_data[24][95] = 0;
        pixel_data[24][96] = 0;
        pixel_data[24][97] = 0;
        pixel_data[24][98] = 0;
        pixel_data[24][99] = 0; // y=24
        pixel_data[25][0] = 0;
        pixel_data[25][1] = 0;
        pixel_data[25][2] = 0;
        pixel_data[25][3] = 0;
        pixel_data[25][4] = 0;
        pixel_data[25][5] = 0;
        pixel_data[25][6] = 0;
        pixel_data[25][7] = 0;
        pixel_data[25][8] = 0;
        pixel_data[25][9] = 0;
        pixel_data[25][10] = 0;
        pixel_data[25][11] = 0;
        pixel_data[25][12] = 0;
        pixel_data[25][13] = 0;
        pixel_data[25][14] = 0;
        pixel_data[25][15] = 0;
        pixel_data[25][16] = 0;
        pixel_data[25][17] = 0;
        pixel_data[25][18] = 0;
        pixel_data[25][19] = 0;
        pixel_data[25][20] = 0;
        pixel_data[25][21] = 0;
        pixel_data[25][22] = 0;
        pixel_data[25][23] = 0;
        pixel_data[25][24] = 0;
        pixel_data[25][25] = 0;
        pixel_data[25][26] = 0;
        pixel_data[25][27] = 0;
        pixel_data[25][28] = 0;
        pixel_data[25][29] = 0;
        pixel_data[25][30] = 0;
        pixel_data[25][31] = 0;
        pixel_data[25][32] = 0;
        pixel_data[25][33] = 0;
        pixel_data[25][34] = 0;
        pixel_data[25][35] = 0;
        pixel_data[25][36] = 0;
        pixel_data[25][37] = 0;
        pixel_data[25][38] = 0;
        pixel_data[25][39] = 0;
        pixel_data[25][40] = 0;
        pixel_data[25][41] = 0;
        pixel_data[25][42] = 0;
        pixel_data[25][43] = 0;
        pixel_data[25][44] = 0;
        pixel_data[25][45] = 0;
        pixel_data[25][46] = 0;
        pixel_data[25][47] = 0;
        pixel_data[25][48] = 0;
        pixel_data[25][49] = 0;
        pixel_data[25][50] = 0;
        pixel_data[25][51] = 0;
        pixel_data[25][52] = 0;
        pixel_data[25][53] = 0;
        pixel_data[25][54] = 0;
        pixel_data[25][55] = 0;
        pixel_data[25][56] = 0;
        pixel_data[25][57] = 0;
        pixel_data[25][58] = 0;
        pixel_data[25][59] = 0;
        pixel_data[25][60] = 0;
        pixel_data[25][61] = 0;
        pixel_data[25][62] = 0;
        pixel_data[25][63] = 0;
        pixel_data[25][64] = 0;
        pixel_data[25][65] = 0;
        pixel_data[25][66] = 0;
        pixel_data[25][67] = 0;
        pixel_data[25][68] = 0;
        pixel_data[25][69] = 0;
        pixel_data[25][70] = 0;
        pixel_data[25][71] = 0;
        pixel_data[25][72] = 0;
        pixel_data[25][73] = 0;
        pixel_data[25][74] = 0;
        pixel_data[25][75] = 0;
        pixel_data[25][76] = 0;
        pixel_data[25][77] = 0;
        pixel_data[25][78] = 0;
        pixel_data[25][79] = 0;
        pixel_data[25][80] = 0;
        pixel_data[25][81] = 0;
        pixel_data[25][82] = 0;
        pixel_data[25][83] = 0;
        pixel_data[25][84] = 0;
        pixel_data[25][85] = 0;
        pixel_data[25][86] = 0;
        pixel_data[25][87] = 0;
        pixel_data[25][88] = 0;
        pixel_data[25][89] = 0;
        pixel_data[25][90] = 0;
        pixel_data[25][91] = 0;
        pixel_data[25][92] = 0;
        pixel_data[25][93] = 0;
        pixel_data[25][94] = 0;
        pixel_data[25][95] = 0;
        pixel_data[25][96] = 0;
        pixel_data[25][97] = 0;
        pixel_data[25][98] = 0;
        pixel_data[25][99] = 0; // y=25
        pixel_data[26][0] = 0;
        pixel_data[26][1] = 0;
        pixel_data[26][2] = 0;
        pixel_data[26][3] = 0;
        pixel_data[26][4] = 0;
        pixel_data[26][5] = 0;
        pixel_data[26][6] = 0;
        pixel_data[26][7] = 0;
        pixel_data[26][8] = 0;
        pixel_data[26][9] = 0;
        pixel_data[26][10] = 0;
        pixel_data[26][11] = 0;
        pixel_data[26][12] = 0;
        pixel_data[26][13] = 0;
        pixel_data[26][14] = 0;
        pixel_data[26][15] = 0;
        pixel_data[26][16] = 0;
        pixel_data[26][17] = 0;
        pixel_data[26][18] = 0;
        pixel_data[26][19] = 0;
        pixel_data[26][20] = 0;
        pixel_data[26][21] = 0;
        pixel_data[26][22] = 0;
        pixel_data[26][23] = 0;
        pixel_data[26][24] = 0;
        pixel_data[26][25] = 0;
        pixel_data[26][26] = 0;
        pixel_data[26][27] = 0;
        pixel_data[26][28] = 0;
        pixel_data[26][29] = 0;
        pixel_data[26][30] = 0;
        pixel_data[26][31] = 0;
        pixel_data[26][32] = 0;
        pixel_data[26][33] = 0;
        pixel_data[26][34] = 0;
        pixel_data[26][35] = 0;
        pixel_data[26][36] = 0;
        pixel_data[26][37] = 0;
        pixel_data[26][38] = 0;
        pixel_data[26][39] = 0;
        pixel_data[26][40] = 0;
        pixel_data[26][41] = 0;
        pixel_data[26][42] = 0;
        pixel_data[26][43] = 0;
        pixel_data[26][44] = 0;
        pixel_data[26][45] = 0;
        pixel_data[26][46] = 0;
        pixel_data[26][47] = 0;
        pixel_data[26][48] = 0;
        pixel_data[26][49] = 0;
        pixel_data[26][50] = 0;
        pixel_data[26][51] = 0;
        pixel_data[26][52] = 0;
        pixel_data[26][53] = 0;
        pixel_data[26][54] = 0;
        pixel_data[26][55] = 0;
        pixel_data[26][56] = 0;
        pixel_data[26][57] = 0;
        pixel_data[26][58] = 0;
        pixel_data[26][59] = 0;
        pixel_data[26][60] = 0;
        pixel_data[26][61] = 0;
        pixel_data[26][62] = 0;
        pixel_data[26][63] = 0;
        pixel_data[26][64] = 0;
        pixel_data[26][65] = 0;
        pixel_data[26][66] = 0;
        pixel_data[26][67] = 0;
        pixel_data[26][68] = 0;
        pixel_data[26][69] = 0;
        pixel_data[26][70] = 0;
        pixel_data[26][71] = 0;
        pixel_data[26][72] = 0;
        pixel_data[26][73] = 0;
        pixel_data[26][74] = 0;
        pixel_data[26][75] = 0;
        pixel_data[26][76] = 0;
        pixel_data[26][77] = 0;
        pixel_data[26][78] = 0;
        pixel_data[26][79] = 0;
        pixel_data[26][80] = 0;
        pixel_data[26][81] = 0;
        pixel_data[26][82] = 0;
        pixel_data[26][83] = 0;
        pixel_data[26][84] = 0;
        pixel_data[26][85] = 0;
        pixel_data[26][86] = 0;
        pixel_data[26][87] = 0;
        pixel_data[26][88] = 0;
        pixel_data[26][89] = 0;
        pixel_data[26][90] = 0;
        pixel_data[26][91] = 0;
        pixel_data[26][92] = 0;
        pixel_data[26][93] = 0;
        pixel_data[26][94] = 0;
        pixel_data[26][95] = 0;
        pixel_data[26][96] = 0;
        pixel_data[26][97] = 0;
        pixel_data[26][98] = 0;
        pixel_data[26][99] = 0; // y=26
        pixel_data[27][0] = 0;
        pixel_data[27][1] = 0;
        pixel_data[27][2] = 0;
        pixel_data[27][3] = 0;
        pixel_data[27][4] = 0;
        pixel_data[27][5] = 0;
        pixel_data[27][6] = 0;
        pixel_data[27][7] = 0;
        pixel_data[27][8] = 0;
        pixel_data[27][9] = 0;
        pixel_data[27][10] = 0;
        pixel_data[27][11] = 0;
        pixel_data[27][12] = 0;
        pixel_data[27][13] = 1;
        pixel_data[27][14] = 1;
        pixel_data[27][15] = 15;
        pixel_data[27][16] = 0;
        pixel_data[27][17] = 0;
        pixel_data[27][18] = 0;
        pixel_data[27][19] = 0;
        pixel_data[27][20] = 0;
        pixel_data[27][21] = 0;
        pixel_data[27][22] = 0;
        pixel_data[27][23] = 0;
        pixel_data[27][24] = 0;
        pixel_data[27][25] = 0;
        pixel_data[27][26] = 0;
        pixel_data[27][27] = 0;
        pixel_data[27][28] = 0;
        pixel_data[27][29] = 0;
        pixel_data[27][30] = 0;
        pixel_data[27][31] = 0;
        pixel_data[27][32] = 0;
        pixel_data[27][33] = 0;
        pixel_data[27][34] = 0;
        pixel_data[27][35] = 0;
        pixel_data[27][36] = 0;
        pixel_data[27][37] = 0;
        pixel_data[27][38] = 0;
        pixel_data[27][39] = 0;
        pixel_data[27][40] = 0;
        pixel_data[27][41] = 0;
        pixel_data[27][42] = 0;
        pixel_data[27][43] = 0;
        pixel_data[27][44] = 0;
        pixel_data[27][45] = 0;
        pixel_data[27][46] = 0;
        pixel_data[27][47] = 0;
        pixel_data[27][48] = 0;
        pixel_data[27][49] = 0;
        pixel_data[27][50] = 0;
        pixel_data[27][51] = 0;
        pixel_data[27][52] = 0;
        pixel_data[27][53] = 0;
        pixel_data[27][54] = 0;
        pixel_data[27][55] = 0;
        pixel_data[27][56] = 0;
        pixel_data[27][57] = 0;
        pixel_data[27][58] = 0;
        pixel_data[27][59] = 0;
        pixel_data[27][60] = 0;
        pixel_data[27][61] = 0;
        pixel_data[27][62] = 0;
        pixel_data[27][63] = 0;
        pixel_data[27][64] = 0;
        pixel_data[27][65] = 0;
        pixel_data[27][66] = 0;
        pixel_data[27][67] = 0;
        pixel_data[27][68] = 0;
        pixel_data[27][69] = 0;
        pixel_data[27][70] = 0;
        pixel_data[27][71] = 0;
        pixel_data[27][72] = 0;
        pixel_data[27][73] = 0;
        pixel_data[27][74] = 0;
        pixel_data[27][75] = 0;
        pixel_data[27][76] = 0;
        pixel_data[27][77] = 0;
        pixel_data[27][78] = 0;
        pixel_data[27][79] = 0;
        pixel_data[27][80] = 0;
        pixel_data[27][81] = 0;
        pixel_data[27][82] = 0;
        pixel_data[27][83] = 0;
        pixel_data[27][84] = 0;
        pixel_data[27][85] = 0;
        pixel_data[27][86] = 0;
        pixel_data[27][87] = 0;
        pixel_data[27][88] = 0;
        pixel_data[27][89] = 0;
        pixel_data[27][90] = 0;
        pixel_data[27][91] = 0;
        pixel_data[27][92] = 0;
        pixel_data[27][93] = 0;
        pixel_data[27][94] = 0;
        pixel_data[27][95] = 0;
        pixel_data[27][96] = 0;
        pixel_data[27][97] = 0;
        pixel_data[27][98] = 0;
        pixel_data[27][99] = 0; // y=27
        pixel_data[28][0] = 0;
        pixel_data[28][1] = 0;
        pixel_data[28][2] = 0;
        pixel_data[28][3] = 0;
        pixel_data[28][4] = 0;
        pixel_data[28][5] = 0;
        pixel_data[28][6] = 0;
        pixel_data[28][7] = 0;
        pixel_data[28][8] = 0;
        pixel_data[28][9] = 0;
        pixel_data[28][10] = 0;
        pixel_data[28][11] = 1;
        pixel_data[28][12] = 7;
        pixel_data[28][13] = 8;
        pixel_data[28][14] = 4;
        pixel_data[28][15] = 6;
        pixel_data[28][16] = 5;
        pixel_data[28][17] = 7;
        pixel_data[28][18] = 1;
        pixel_data[28][19] = 0;
        pixel_data[28][20] = 0;
        pixel_data[28][21] = 0;
        pixel_data[28][22] = 0;
        pixel_data[28][23] = 0;
        pixel_data[28][24] = 0;
        pixel_data[28][25] = 0;
        pixel_data[28][26] = 0;
        pixel_data[28][27] = 0;
        pixel_data[28][28] = 0;
        pixel_data[28][29] = 0;
        pixel_data[28][30] = 0;
        pixel_data[28][31] = 0;
        pixel_data[28][32] = 0;
        pixel_data[28][33] = 0;
        pixel_data[28][34] = 0;
        pixel_data[28][35] = 0;
        pixel_data[28][36] = 0;
        pixel_data[28][37] = 0;
        pixel_data[28][38] = 0;
        pixel_data[28][39] = 0;
        pixel_data[28][40] = 0;
        pixel_data[28][41] = 0;
        pixel_data[28][42] = 0;
        pixel_data[28][43] = 0;
        pixel_data[28][44] = 0;
        pixel_data[28][45] = 0;
        pixel_data[28][46] = 0;
        pixel_data[28][47] = 0;
        pixel_data[28][48] = 0;
        pixel_data[28][49] = 0;
        pixel_data[28][50] = 0;
        pixel_data[28][51] = 0;
        pixel_data[28][52] = 0;
        pixel_data[28][53] = 0;
        pixel_data[28][54] = 0;
        pixel_data[28][55] = 0;
        pixel_data[28][56] = 0;
        pixel_data[28][57] = 0;
        pixel_data[28][58] = 0;
        pixel_data[28][59] = 0;
        pixel_data[28][60] = 0;
        pixel_data[28][61] = 0;
        pixel_data[28][62] = 0;
        pixel_data[28][63] = 0;
        pixel_data[28][64] = 0;
        pixel_data[28][65] = 0;
        pixel_data[28][66] = 0;
        pixel_data[28][67] = 0;
        pixel_data[28][68] = 0;
        pixel_data[28][69] = 0;
        pixel_data[28][70] = 0;
        pixel_data[28][71] = 0;
        pixel_data[28][72] = 0;
        pixel_data[28][73] = 0;
        pixel_data[28][74] = 0;
        pixel_data[28][75] = 0;
        pixel_data[28][76] = 0;
        pixel_data[28][77] = 0;
        pixel_data[28][78] = 0;
        pixel_data[28][79] = 0;
        pixel_data[28][80] = 0;
        pixel_data[28][81] = 0;
        pixel_data[28][82] = 0;
        pixel_data[28][83] = 0;
        pixel_data[28][84] = 0;
        pixel_data[28][85] = 0;
        pixel_data[28][86] = 0;
        pixel_data[28][87] = 0;
        pixel_data[28][88] = 0;
        pixel_data[28][89] = 0;
        pixel_data[28][90] = 0;
        pixel_data[28][91] = 0;
        pixel_data[28][92] = 0;
        pixel_data[28][93] = 0;
        pixel_data[28][94] = 0;
        pixel_data[28][95] = 0;
        pixel_data[28][96] = 0;
        pixel_data[28][97] = 0;
        pixel_data[28][98] = 0;
        pixel_data[28][99] = 0; // y=28
        pixel_data[29][0] = 0;
        pixel_data[29][1] = 0;
        pixel_data[29][2] = 0;
        pixel_data[29][3] = 0;
        pixel_data[29][4] = 0;
        pixel_data[29][5] = 0;
        pixel_data[29][6] = 0;
        pixel_data[29][7] = 0;
        pixel_data[29][8] = 0;
        pixel_data[29][9] = 0;
        pixel_data[29][10] = 2;
        pixel_data[29][11] = 8;
        pixel_data[29][12] = 6;
        pixel_data[29][13] = 6;
        pixel_data[29][14] = 6;
        pixel_data[29][15] = 6;
        pixel_data[29][16] = 6;
        pixel_data[29][17] = 6;
        pixel_data[29][18] = 6;
        pixel_data[29][19] = 6;
        pixel_data[29][20] = 11;
        pixel_data[29][21] = 15;
        pixel_data[29][22] = 0;
        pixel_data[29][23] = 0;
        pixel_data[29][24] = 0;
        pixel_data[29][25] = 0;
        pixel_data[29][26] = 0;
        pixel_data[29][27] = 0;
        pixel_data[29][28] = 0;
        pixel_data[29][29] = 0;
        pixel_data[29][30] = 0;
        pixel_data[29][31] = 1;
        pixel_data[29][32] = 15;
        pixel_data[29][33] = 15;
        pixel_data[29][34] = 15;
        pixel_data[29][35] = 1;
        pixel_data[29][36] = 0;
        pixel_data[29][37] = 0;
        pixel_data[29][38] = 0;
        pixel_data[29][39] = 0;
        pixel_data[29][40] = 0;
        pixel_data[29][41] = 0;
        pixel_data[29][42] = 0;
        pixel_data[29][43] = 0;
        pixel_data[29][44] = 0;
        pixel_data[29][45] = 0;
        pixel_data[29][46] = 0;
        pixel_data[29][47] = 0;
        pixel_data[29][48] = 0;
        pixel_data[29][49] = 0;
        pixel_data[29][50] = 0;
        pixel_data[29][51] = 0;
        pixel_data[29][52] = 0;
        pixel_data[29][53] = 0;
        pixel_data[29][54] = 0;
        pixel_data[29][55] = 0;
        pixel_data[29][56] = 0;
        pixel_data[29][57] = 0;
        pixel_data[29][58] = 0;
        pixel_data[29][59] = 0;
        pixel_data[29][60] = 0;
        pixel_data[29][61] = 0;
        pixel_data[29][62] = 0;
        pixel_data[29][63] = 0;
        pixel_data[29][64] = 0;
        pixel_data[29][65] = 0;
        pixel_data[29][66] = 0;
        pixel_data[29][67] = 0;
        pixel_data[29][68] = 0;
        pixel_data[29][69] = 0;
        pixel_data[29][70] = 0;
        pixel_data[29][71] = 0;
        pixel_data[29][72] = 0;
        pixel_data[29][73] = 0;
        pixel_data[29][74] = 0;
        pixel_data[29][75] = 0;
        pixel_data[29][76] = 0;
        pixel_data[29][77] = 0;
        pixel_data[29][78] = 0;
        pixel_data[29][79] = 0;
        pixel_data[29][80] = 0;
        pixel_data[29][81] = 0;
        pixel_data[29][82] = 0;
        pixel_data[29][83] = 0;
        pixel_data[29][84] = 0;
        pixel_data[29][85] = 0;
        pixel_data[29][86] = 0;
        pixel_data[29][87] = 0;
        pixel_data[29][88] = 0;
        pixel_data[29][89] = 0;
        pixel_data[29][90] = 0;
        pixel_data[29][91] = 0;
        pixel_data[29][92] = 0;
        pixel_data[29][93] = 0;
        pixel_data[29][94] = 0;
        pixel_data[29][95] = 0;
        pixel_data[29][96] = 0;
        pixel_data[29][97] = 0;
        pixel_data[29][98] = 0;
        pixel_data[29][99] = 0; // y=29
        pixel_data[30][0] = 0;
        pixel_data[30][1] = 0;
        pixel_data[30][2] = 0;
        pixel_data[30][3] = 0;
        pixel_data[30][4] = 0;
        pixel_data[30][5] = 0;
        pixel_data[30][6] = 0;
        pixel_data[30][7] = 0;
        pixel_data[30][8] = 0;
        pixel_data[30][9] = 0;
        pixel_data[30][10] = 7;
        pixel_data[30][11] = 6;
        pixel_data[30][12] = 6;
        pixel_data[30][13] = 6;
        pixel_data[30][14] = 6;
        pixel_data[30][15] = 6;
        pixel_data[30][16] = 6;
        pixel_data[30][17] = 6;
        pixel_data[30][18] = 6;
        pixel_data[30][19] = 6;
        pixel_data[30][20] = 6;
        pixel_data[30][21] = 8;
        pixel_data[30][22] = 6;
        pixel_data[30][23] = 4;
        pixel_data[30][24] = 5;
        pixel_data[30][25] = 5;
        pixel_data[30][26] = 7;
        pixel_data[30][27] = 12;
        pixel_data[30][28] = 2;
        pixel_data[30][29] = 2;
        pixel_data[30][30] = 2;
        pixel_data[30][31] = 11;
        pixel_data[30][32] = 10;
        pixel_data[30][33] = 7;
        pixel_data[30][34] = 7;
        pixel_data[30][35] = 7;
        pixel_data[30][36] = 7;
        pixel_data[30][37] = 12;
        pixel_data[30][38] = 14;
        pixel_data[30][39] = 0;
        pixel_data[30][40] = 0;
        pixel_data[30][41] = 0;
        pixel_data[30][42] = 0;
        pixel_data[30][43] = 0;
        pixel_data[30][44] = 0;
        pixel_data[30][45] = 0;
        pixel_data[30][46] = 0;
        pixel_data[30][47] = 0;
        pixel_data[30][48] = 0;
        pixel_data[30][49] = 0;
        pixel_data[30][50] = 0;
        pixel_data[30][51] = 0;
        pixel_data[30][52] = 0;
        pixel_data[30][53] = 0;
        pixel_data[30][54] = 0;
        pixel_data[30][55] = 0;
        pixel_data[30][56] = 0;
        pixel_data[30][57] = 0;
        pixel_data[30][58] = 0;
        pixel_data[30][59] = 0;
        pixel_data[30][60] = 0;
        pixel_data[30][61] = 0;
        pixel_data[30][62] = 0;
        pixel_data[30][63] = 0;
        pixel_data[30][64] = 0;
        pixel_data[30][65] = 0;
        pixel_data[30][66] = 0;
        pixel_data[30][67] = 0;
        pixel_data[30][68] = 0;
        pixel_data[30][69] = 0;
        pixel_data[30][70] = 0;
        pixel_data[30][71] = 0;
        pixel_data[30][72] = 0;
        pixel_data[30][73] = 0;
        pixel_data[30][74] = 0;
        pixel_data[30][75] = 0;
        pixel_data[30][76] = 0;
        pixel_data[30][77] = 0;
        pixel_data[30][78] = 0;
        pixel_data[30][79] = 0;
        pixel_data[30][80] = 0;
        pixel_data[30][81] = 0;
        pixel_data[30][82] = 0;
        pixel_data[30][83] = 0;
        pixel_data[30][84] = 0;
        pixel_data[30][85] = 0;
        pixel_data[30][86] = 0;
        pixel_data[30][87] = 0;
        pixel_data[30][88] = 0;
        pixel_data[30][89] = 0;
        pixel_data[30][90] = 0;
        pixel_data[30][91] = 0;
        pixel_data[30][92] = 0;
        pixel_data[30][93] = 0;
        pixel_data[30][94] = 0;
        pixel_data[30][95] = 0;
        pixel_data[30][96] = 0;
        pixel_data[30][97] = 0;
        pixel_data[30][98] = 0;
        pixel_data[30][99] = 0; // y=30
        pixel_data[31][0] = 0;
        pixel_data[31][1] = 0;
        pixel_data[31][2] = 0;
        pixel_data[31][3] = 0;
        pixel_data[31][4] = 0;
        pixel_data[31][5] = 0;
        pixel_data[31][6] = 0;
        pixel_data[31][7] = 0;
        pixel_data[31][8] = 0;
        pixel_data[31][9] = 7;
        pixel_data[31][10] = 8;
        pixel_data[31][11] = 6;
        pixel_data[31][12] = 6;
        pixel_data[31][13] = 6;
        pixel_data[31][14] = 6;
        pixel_data[31][15] = 6;
        pixel_data[31][16] = 6;
        pixel_data[31][17] = 6;
        pixel_data[31][18] = 6;
        pixel_data[31][19] = 6;
        pixel_data[31][20] = 6;
        pixel_data[31][21] = 6;
        pixel_data[31][22] = 6;
        pixel_data[31][23] = 6;
        pixel_data[31][24] = 6;
        pixel_data[31][25] = 8;
        pixel_data[31][26] = 9;
        pixel_data[31][27] = 9;
        pixel_data[31][28] = 9;
        pixel_data[31][29] = 9;
        pixel_data[31][30] = 10;
        pixel_data[31][31] = 10;
        pixel_data[31][32] = 10;
        pixel_data[31][33] = 10;
        pixel_data[31][34] = 10;
        pixel_data[31][35] = 9;
        pixel_data[31][36] = 9;
        pixel_data[31][37] = 10;
        pixel_data[31][38] = 11;
        pixel_data[31][39] = 5;
        pixel_data[31][40] = 2;
        pixel_data[31][41] = 7;
        pixel_data[31][42] = 1;
        pixel_data[31][43] = 0;
        pixel_data[31][44] = 0;
        pixel_data[31][45] = 0;
        pixel_data[31][46] = 0;
        pixel_data[31][47] = 0;
        pixel_data[31][48] = 0;
        pixel_data[31][49] = 0;
        pixel_data[31][50] = 0;
        pixel_data[31][51] = 0;
        pixel_data[31][52] = 0;
        pixel_data[31][53] = 0;
        pixel_data[31][54] = 0;
        pixel_data[31][55] = 0;
        pixel_data[31][56] = 0;
        pixel_data[31][57] = 0;
        pixel_data[31][58] = 0;
        pixel_data[31][59] = 0;
        pixel_data[31][60] = 0;
        pixel_data[31][61] = 0;
        pixel_data[31][62] = 0;
        pixel_data[31][63] = 0;
        pixel_data[31][64] = 0;
        pixel_data[31][65] = 0;
        pixel_data[31][66] = 0;
        pixel_data[31][67] = 0;
        pixel_data[31][68] = 0;
        pixel_data[31][69] = 0;
        pixel_data[31][70] = 0;
        pixel_data[31][71] = 0;
        pixel_data[31][72] = 0;
        pixel_data[31][73] = 0;
        pixel_data[31][74] = 0;
        pixel_data[31][75] = 0;
        pixel_data[31][76] = 0;
        pixel_data[31][77] = 0;
        pixel_data[31][78] = 0;
        pixel_data[31][79] = 0;
        pixel_data[31][80] = 0;
        pixel_data[31][81] = 0;
        pixel_data[31][82] = 0;
        pixel_data[31][83] = 0;
        pixel_data[31][84] = 0;
        pixel_data[31][85] = 0;
        pixel_data[31][86] = 0;
        pixel_data[31][87] = 0;
        pixel_data[31][88] = 0;
        pixel_data[31][89] = 0;
        pixel_data[31][90] = 0;
        pixel_data[31][91] = 0;
        pixel_data[31][92] = 0;
        pixel_data[31][93] = 0;
        pixel_data[31][94] = 0;
        pixel_data[31][95] = 0;
        pixel_data[31][96] = 0;
        pixel_data[31][97] = 0;
        pixel_data[31][98] = 0;
        pixel_data[31][99] = 0; // y=31
        pixel_data[32][0] = 0;
        pixel_data[32][1] = 0;
        pixel_data[32][2] = 0;
        pixel_data[32][3] = 0;
        pixel_data[32][4] = 0;
        pixel_data[32][5] = 0;
        pixel_data[32][6] = 0;
        pixel_data[32][7] = 0;
        pixel_data[32][8] = 0;
        pixel_data[32][9] = 5;
        pixel_data[32][10] = 6;
        pixel_data[32][11] = 6;
        pixel_data[32][12] = 6;
        pixel_data[32][13] = 6;
        pixel_data[32][14] = 6;
        pixel_data[32][15] = 6;
        pixel_data[32][16] = 6;
        pixel_data[32][17] = 6;
        pixel_data[32][18] = 6;
        pixel_data[32][19] = 6;
        pixel_data[32][20] = 6;
        pixel_data[32][21] = 6;
        pixel_data[32][22] = 6;
        pixel_data[32][23] = 8;
        pixel_data[32][24] = 8;
        pixel_data[32][25] = 9;
        pixel_data[32][26] = 9;
        pixel_data[32][27] = 9;
        pixel_data[32][28] = 10;
        pixel_data[32][29] = 9;
        pixel_data[32][30] = 10;
        pixel_data[32][31] = 10;
        pixel_data[32][32] = 10;
        pixel_data[32][33] = 10;
        pixel_data[32][34] = 10;
        pixel_data[32][35] = 10;
        pixel_data[32][36] = 10;
        pixel_data[32][37] = 9;
        pixel_data[32][38] = 9;
        pixel_data[32][39] = 10;
        pixel_data[32][40] = 7;
        pixel_data[32][41] = 10;
        pixel_data[32][42] = 5;
        pixel_data[32][43] = 11;
        pixel_data[32][44] = 12;
        pixel_data[32][45] = 1;
        pixel_data[32][46] = 0;
        pixel_data[32][47] = 0;
        pixel_data[32][48] = 0;
        pixel_data[32][49] = 0;
        pixel_data[32][50] = 0;
        pixel_data[32][51] = 0;
        pixel_data[32][52] = 0;
        pixel_data[32][53] = 0;
        pixel_data[32][54] = 0;
        pixel_data[32][55] = 0;
        pixel_data[32][56] = 0;
        pixel_data[32][57] = 0;
        pixel_data[32][58] = 0;
        pixel_data[32][59] = 0;
        pixel_data[32][60] = 0;
        pixel_data[32][61] = 0;
        pixel_data[32][62] = 0;
        pixel_data[32][63] = 0;
        pixel_data[32][64] = 0;
        pixel_data[32][65] = 0;
        pixel_data[32][66] = 0;
        pixel_data[32][67] = 0;
        pixel_data[32][68] = 0;
        pixel_data[32][69] = 0;
        pixel_data[32][70] = 0;
        pixel_data[32][71] = 0;
        pixel_data[32][72] = 0;
        pixel_data[32][73] = 0;
        pixel_data[32][74] = 0;
        pixel_data[32][75] = 0;
        pixel_data[32][76] = 0;
        pixel_data[32][77] = 0;
        pixel_data[32][78] = 0;
        pixel_data[32][79] = 0;
        pixel_data[32][80] = 0;
        pixel_data[32][81] = 0;
        pixel_data[32][82] = 0;
        pixel_data[32][83] = 0;
        pixel_data[32][84] = 0;
        pixel_data[32][85] = 0;
        pixel_data[32][86] = 0;
        pixel_data[32][87] = 0;
        pixel_data[32][88] = 0;
        pixel_data[32][89] = 0;
        pixel_data[32][90] = 0;
        pixel_data[32][91] = 0;
        pixel_data[32][92] = 0;
        pixel_data[32][93] = 0;
        pixel_data[32][94] = 0;
        pixel_data[32][95] = 0;
        pixel_data[32][96] = 0;
        pixel_data[32][97] = 0;
        pixel_data[32][98] = 0;
        pixel_data[32][99] = 0; // y=32
        pixel_data[33][0] = 0;
        pixel_data[33][1] = 0;
        pixel_data[33][2] = 0;
        pixel_data[33][3] = 0;
        pixel_data[33][4] = 0;
        pixel_data[33][5] = 0;
        pixel_data[33][6] = 0;
        pixel_data[33][7] = 0;
        pixel_data[33][8] = 0;
        pixel_data[33][9] = 5;
        pixel_data[33][10] = 6;
        pixel_data[33][11] = 6;
        pixel_data[33][12] = 6;
        pixel_data[33][13] = 6;
        pixel_data[33][14] = 6;
        pixel_data[33][15] = 6;
        pixel_data[33][16] = 6;
        pixel_data[33][17] = 6;
        pixel_data[33][18] = 6;
        pixel_data[33][19] = 6;
        pixel_data[33][20] = 8;
        pixel_data[33][21] = 8;
        pixel_data[33][22] = 8;
        pixel_data[33][23] = 9;
        pixel_data[33][24] = 9;
        pixel_data[33][25] = 9;
        pixel_data[33][26] = 10;
        pixel_data[33][27] = 10;
        pixel_data[33][28] = 10;
        pixel_data[33][29] = 10;
        pixel_data[33][30] = 10;
        pixel_data[33][31] = 11;
        pixel_data[33][32] = 10;
        pixel_data[33][33] = 10;
        pixel_data[33][34] = 10;
        pixel_data[33][35] = 10;
        pixel_data[33][36] = 10;
        pixel_data[33][37] = 10;
        pixel_data[33][38] = 10;
        pixel_data[33][39] = 10;
        pixel_data[33][40] = 9;
        pixel_data[33][41] = 9;
        pixel_data[33][42] = 9;
        pixel_data[33][43] = 10;
        pixel_data[33][44] = 9;
        pixel_data[33][45] = 7;
        pixel_data[33][46] = 10;
        pixel_data[33][47] = 11;
        pixel_data[33][48] = 2;
        pixel_data[33][49] = 1;
        pixel_data[33][50] = 1;
        pixel_data[33][51] = 0;
        pixel_data[33][52] = 0;
        pixel_data[33][53] = 0;
        pixel_data[33][54] = 0;
        pixel_data[33][55] = 0;
        pixel_data[33][56] = 0;
        pixel_data[33][57] = 0;
        pixel_data[33][58] = 0;
        pixel_data[33][59] = 0;
        pixel_data[33][60] = 0;
        pixel_data[33][61] = 0;
        pixel_data[33][62] = 0;
        pixel_data[33][63] = 0;
        pixel_data[33][64] = 0;
        pixel_data[33][65] = 0;
        pixel_data[33][66] = 0;
        pixel_data[33][67] = 0;
        pixel_data[33][68] = 0;
        pixel_data[33][69] = 0;
        pixel_data[33][70] = 0;
        pixel_data[33][71] = 0;
        pixel_data[33][72] = 0;
        pixel_data[33][73] = 0;
        pixel_data[33][74] = 0;
        pixel_data[33][75] = 0;
        pixel_data[33][76] = 0;
        pixel_data[33][77] = 0;
        pixel_data[33][78] = 0;
        pixel_data[33][79] = 0;
        pixel_data[33][80] = 0;
        pixel_data[33][81] = 0;
        pixel_data[33][82] = 0;
        pixel_data[33][83] = 0;
        pixel_data[33][84] = 0;
        pixel_data[33][85] = 0;
        pixel_data[33][86] = 0;
        pixel_data[33][87] = 0;
        pixel_data[33][88] = 0;
        pixel_data[33][89] = 0;
        pixel_data[33][90] = 0;
        pixel_data[33][91] = 0;
        pixel_data[33][92] = 0;
        pixel_data[33][93] = 0;
        pixel_data[33][94] = 0;
        pixel_data[33][95] = 0;
        pixel_data[33][96] = 0;
        pixel_data[33][97] = 0;
        pixel_data[33][98] = 0;
        pixel_data[33][99] = 0; // y=33
        pixel_data[34][0] = 0;
        pixel_data[34][1] = 0;
        pixel_data[34][2] = 0;
        pixel_data[34][3] = 0;
        pixel_data[34][4] = 0;
        pixel_data[34][5] = 0;
        pixel_data[34][6] = 0;
        pixel_data[34][7] = 0;
        pixel_data[34][8] = 0;
        pixel_data[34][9] = 2;
        pixel_data[34][10] = 6;
        pixel_data[34][11] = 6;
        pixel_data[34][12] = 6;
        pixel_data[34][13] = 6;
        pixel_data[34][14] = 6;
        pixel_data[34][15] = 6;
        pixel_data[34][16] = 6;
        pixel_data[34][17] = 6;
        pixel_data[34][18] = 6;
        pixel_data[34][19] = 8;
        pixel_data[34][20] = 8;
        pixel_data[34][21] = 8;
        pixel_data[34][22] = 9;
        pixel_data[34][23] = 9;
        pixel_data[34][24] = 10;
        pixel_data[34][25] = 10;
        pixel_data[34][26] = 10;
        pixel_data[34][27] = 10;
        pixel_data[34][28] = 11;
        pixel_data[34][29] = 11;
        pixel_data[34][30] = 11;
        pixel_data[34][31] = 11;
        pixel_data[34][32] = 11;
        pixel_data[34][33] = 11;
        pixel_data[34][34] = 11;
        pixel_data[34][35] = 11;
        pixel_data[34][36] = 11;
        pixel_data[34][37] = 10;
        pixel_data[34][38] = 10;
        pixel_data[34][39] = 10;
        pixel_data[34][40] = 9;
        pixel_data[34][41] = 10;
        pixel_data[34][42] = 10;
        pixel_data[34][43] = 10;
        pixel_data[34][44] = 10;
        pixel_data[34][45] = 10;
        pixel_data[34][46] = 10;
        pixel_data[34][47] = 10;
        pixel_data[34][48] = 10;
        pixel_data[34][49] = 10;
        pixel_data[34][50] = 7;
        pixel_data[34][51] = 12;
        pixel_data[34][52] = 14;
        pixel_data[34][53] = 1;
        pixel_data[34][54] = 0;
        pixel_data[34][55] = 0;
        pixel_data[34][56] = 0;
        pixel_data[34][57] = 0;
        pixel_data[34][58] = 0;
        pixel_data[34][59] = 0;
        pixel_data[34][60] = 0;
        pixel_data[34][61] = 0;
        pixel_data[34][62] = 0;
        pixel_data[34][63] = 0;
        pixel_data[34][64] = 0;
        pixel_data[34][65] = 0;
        pixel_data[34][66] = 0;
        pixel_data[34][67] = 0;
        pixel_data[34][68] = 0;
        pixel_data[34][69] = 0;
        pixel_data[34][70] = 0;
        pixel_data[34][71] = 0;
        pixel_data[34][72] = 0;
        pixel_data[34][73] = 0;
        pixel_data[34][74] = 0;
        pixel_data[34][75] = 0;
        pixel_data[34][76] = 0;
        pixel_data[34][77] = 0;
        pixel_data[34][78] = 0;
        pixel_data[34][79] = 0;
        pixel_data[34][80] = 0;
        pixel_data[34][81] = 0;
        pixel_data[34][82] = 0;
        pixel_data[34][83] = 0;
        pixel_data[34][84] = 0;
        pixel_data[34][85] = 0;
        pixel_data[34][86] = 0;
        pixel_data[34][87] = 0;
        pixel_data[34][88] = 0;
        pixel_data[34][89] = 0;
        pixel_data[34][90] = 0;
        pixel_data[34][91] = 0;
        pixel_data[34][92] = 0;
        pixel_data[34][93] = 0;
        pixel_data[34][94] = 0;
        pixel_data[34][95] = 0;
        pixel_data[34][96] = 0;
        pixel_data[34][97] = 0;
        pixel_data[34][98] = 0;
        pixel_data[34][99] = 0; // y=34
        pixel_data[35][0] = 0;
        pixel_data[35][1] = 0;
        pixel_data[35][2] = 0;
        pixel_data[35][3] = 0;
        pixel_data[35][4] = 0;
        pixel_data[35][5] = 0;
        pixel_data[35][6] = 0;
        pixel_data[35][7] = 0;
        pixel_data[35][8] = 0;
        pixel_data[35][9] = 1;
        pixel_data[35][10] = 7;
        pixel_data[35][11] = 6;
        pixel_data[35][12] = 6;
        pixel_data[35][13] = 6;
        pixel_data[35][14] = 6;
        pixel_data[35][15] = 6;
        pixel_data[35][16] = 6;
        pixel_data[35][17] = 6;
        pixel_data[35][18] = 8;
        pixel_data[35][19] = 8;
        pixel_data[35][20] = 8;
        pixel_data[35][21] = 9;
        pixel_data[35][22] = 9;
        pixel_data[35][23] = 10;
        pixel_data[35][24] = 10;
        pixel_data[35][25] = 10;
        pixel_data[35][26] = 10;
        pixel_data[35][27] = 10;
        pixel_data[35][28] = 10;
        pixel_data[35][29] = 11;
        pixel_data[35][30] = 11;
        pixel_data[35][31] = 11;
        pixel_data[35][32] = 11;
        pixel_data[35][33] = 11;
        pixel_data[35][34] = 11;
        pixel_data[35][35] = 11;
        pixel_data[35][36] = 11;
        pixel_data[35][37] = 11;
        pixel_data[35][38] = 10;
        pixel_data[35][39] = 8;
        pixel_data[35][40] = 6;
        pixel_data[35][41] = 6;
        pixel_data[35][42] = 6;
        pixel_data[35][43] = 8;
        pixel_data[35][44] = 8;
        pixel_data[35][45] = 8;
        pixel_data[35][46] = 9;
        pixel_data[35][47] = 10;
        pixel_data[35][48] = 10;
        pixel_data[35][49] = 10;
        pixel_data[35][50] = 11;
        pixel_data[35][51] = 11;
        pixel_data[35][52] = 10;
        pixel_data[35][53] = 12;
        pixel_data[35][54] = 11;
        pixel_data[35][55] = 1;
        pixel_data[35][56] = 0;
        pixel_data[35][57] = 0;
        pixel_data[35][58] = 0;
        pixel_data[35][59] = 0;
        pixel_data[35][60] = 0;
        pixel_data[35][61] = 0;
        pixel_data[35][62] = 0;
        pixel_data[35][63] = 0;
        pixel_data[35][64] = 0;
        pixel_data[35][65] = 0;
        pixel_data[35][66] = 0;
        pixel_data[35][67] = 0;
        pixel_data[35][68] = 0;
        pixel_data[35][69] = 0;
        pixel_data[35][70] = 0;
        pixel_data[35][71] = 0;
        pixel_data[35][72] = 0;
        pixel_data[35][73] = 0;
        pixel_data[35][74] = 0;
        pixel_data[35][75] = 0;
        pixel_data[35][76] = 0;
        pixel_data[35][77] = 0;
        pixel_data[35][78] = 0;
        pixel_data[35][79] = 0;
        pixel_data[35][80] = 0;
        pixel_data[35][81] = 0;
        pixel_data[35][82] = 0;
        pixel_data[35][83] = 0;
        pixel_data[35][84] = 0;
        pixel_data[35][85] = 0;
        pixel_data[35][86] = 0;
        pixel_data[35][87] = 0;
        pixel_data[35][88] = 0;
        pixel_data[35][89] = 0;
        pixel_data[35][90] = 0;
        pixel_data[35][91] = 0;
        pixel_data[35][92] = 0;
        pixel_data[35][93] = 0;
        pixel_data[35][94] = 0;
        pixel_data[35][95] = 0;
        pixel_data[35][96] = 0;
        pixel_data[35][97] = 0;
        pixel_data[35][98] = 0;
        pixel_data[35][99] = 0; // y=35
        pixel_data[36][0] = 0;
        pixel_data[36][1] = 0;
        pixel_data[36][2] = 0;
        pixel_data[36][3] = 0;
        pixel_data[36][4] = 0;
        pixel_data[36][5] = 0;
        pixel_data[36][6] = 0;
        pixel_data[36][7] = 0;
        pixel_data[36][8] = 0;
        pixel_data[36][9] = 0;
        pixel_data[36][10] = 12;
        pixel_data[36][11] = 5;
        pixel_data[36][12] = 6;
        pixel_data[36][13] = 6;
        pixel_data[36][14] = 6;
        pixel_data[36][15] = 6;
        pixel_data[36][16] = 6;
        pixel_data[36][17] = 8;
        pixel_data[36][18] = 8;
        pixel_data[36][19] = 8;
        pixel_data[36][20] = 8;
        pixel_data[36][21] = 9;
        pixel_data[36][22] = 9;
        pixel_data[36][23] = 10;
        pixel_data[36][24] = 10;
        pixel_data[36][25] = 10;
        pixel_data[36][26] = 10;
        pixel_data[36][27] = 10;
        pixel_data[36][28] = 11;
        pixel_data[36][29] = 11;
        pixel_data[36][30] = 11;
        pixel_data[36][31] = 10;
        pixel_data[36][32] = 10;
        pixel_data[36][33] = 10;
        pixel_data[36][34] = 10;
        pixel_data[36][35] = 10;
        pixel_data[36][36] = 10;
        pixel_data[36][37] = 9;
        pixel_data[36][38] = 6;
        pixel_data[36][39] = 4;
        pixel_data[36][40] = 3;
        pixel_data[36][41] = 3;
        pixel_data[36][42] = 3;
        pixel_data[36][43] = 3;
        pixel_data[36][44] = 3;
        pixel_data[36][45] = 3;
        pixel_data[36][46] = 3;
        pixel_data[36][47] = 4;
        pixel_data[36][48] = 6;
        pixel_data[36][49] = 6;
        pixel_data[36][50] = 8;
        pixel_data[36][51] = 10;
        pixel_data[36][52] = 10;
        pixel_data[36][53] = 11;
        pixel_data[36][54] = 11;
        pixel_data[36][55] = 10;
        pixel_data[36][56] = 7;
        pixel_data[36][57] = 7;
        pixel_data[36][58] = 15;
        pixel_data[36][59] = 15;
        pixel_data[36][60] = 0;
        pixel_data[36][61] = 0;
        pixel_data[36][62] = 0;
        pixel_data[36][63] = 0;
        pixel_data[36][64] = 0;
        pixel_data[36][65] = 0;
        pixel_data[36][66] = 0;
        pixel_data[36][67] = 0;
        pixel_data[36][68] = 0;
        pixel_data[36][69] = 0;
        pixel_data[36][70] = 0;
        pixel_data[36][71] = 0;
        pixel_data[36][72] = 0;
        pixel_data[36][73] = 0;
        pixel_data[36][74] = 0;
        pixel_data[36][75] = 0;
        pixel_data[36][76] = 0;
        pixel_data[36][77] = 0;
        pixel_data[36][78] = 0;
        pixel_data[36][79] = 0;
        pixel_data[36][80] = 0;
        pixel_data[36][81] = 0;
        pixel_data[36][82] = 0;
        pixel_data[36][83] = 0;
        pixel_data[36][84] = 0;
        pixel_data[36][85] = 0;
        pixel_data[36][86] = 0;
        pixel_data[36][87] = 0;
        pixel_data[36][88] = 0;
        pixel_data[36][89] = 0;
        pixel_data[36][90] = 0;
        pixel_data[36][91] = 0;
        pixel_data[36][92] = 0;
        pixel_data[36][93] = 0;
        pixel_data[36][94] = 0;
        pixel_data[36][95] = 0;
        pixel_data[36][96] = 0;
        pixel_data[36][97] = 0;
        pixel_data[36][98] = 0;
        pixel_data[36][99] = 0; // y=36
        pixel_data[37][0] = 0;
        pixel_data[37][1] = 0;
        pixel_data[37][2] = 0;
        pixel_data[37][3] = 0;
        pixel_data[37][4] = 0;
        pixel_data[37][5] = 0;
        pixel_data[37][6] = 0;
        pixel_data[37][7] = 0;
        pixel_data[37][8] = 0;
        pixel_data[37][9] = 0;
        pixel_data[37][10] = 0;
        pixel_data[37][11] = 0;
        pixel_data[37][12] = 5;
        pixel_data[37][13] = 8;
        pixel_data[37][14] = 6;
        pixel_data[37][15] = 6;
        pixel_data[37][16] = 6;
        pixel_data[37][17] = 6;
        pixel_data[37][18] = 8;
        pixel_data[37][19] = 8;
        pixel_data[37][20] = 8;
        pixel_data[37][21] = 9;
        pixel_data[37][22] = 9;
        pixel_data[37][23] = 9;
        pixel_data[37][24] = 10;
        pixel_data[37][25] = 10;
        pixel_data[37][26] = 10;
        pixel_data[37][27] = 10;
        pixel_data[37][28] = 11;
        pixel_data[37][29] = 11;
        pixel_data[37][30] = 10;
        pixel_data[37][31] = 10;
        pixel_data[37][32] = 10;
        pixel_data[37][33] = 10;
        pixel_data[37][34] = 10;
        pixel_data[37][35] = 10;
        pixel_data[37][36] = 9;
        pixel_data[37][37] = 8;
        pixel_data[37][38] = 6;
        pixel_data[37][39] = 4;
        pixel_data[37][40] = 4;
        pixel_data[37][41] = 4;
        pixel_data[37][42] = 4;
        pixel_data[37][43] = 3;
        pixel_data[37][44] = 3;
        pixel_data[37][45] = 3;
        pixel_data[37][46] = 3;
        pixel_data[37][47] = 3;
        pixel_data[37][48] = 3;
        pixel_data[37][49] = 3;
        pixel_data[37][50] = 3;
        pixel_data[37][51] = 3;
        pixel_data[37][52] = 4;
        pixel_data[37][53] = 6;
        pixel_data[37][54] = 6;
        pixel_data[37][55] = 6;
        pixel_data[37][56] = 8;
        pixel_data[37][57] = 8;
        pixel_data[37][58] = 6;
        pixel_data[37][59] = 2;
        pixel_data[37][60] = 15;
        pixel_data[37][61] = 7;
        pixel_data[37][62] = 15;
        pixel_data[37][63] = 15;
        pixel_data[37][64] = 0;
        pixel_data[37][65] = 0;
        pixel_data[37][66] = 0;
        pixel_data[37][67] = 0;
        pixel_data[37][68] = 0;
        pixel_data[37][69] = 0;
        pixel_data[37][70] = 0;
        pixel_data[37][71] = 0;
        pixel_data[37][72] = 0;
        pixel_data[37][73] = 0;
        pixel_data[37][74] = 0;
        pixel_data[37][75] = 0;
        pixel_data[37][76] = 0;
        pixel_data[37][77] = 0;
        pixel_data[37][78] = 0;
        pixel_data[37][79] = 0;
        pixel_data[37][80] = 0;
        pixel_data[37][81] = 0;
        pixel_data[37][82] = 0;
        pixel_data[37][83] = 0;
        pixel_data[37][84] = 0;
        pixel_data[37][85] = 0;
        pixel_data[37][86] = 0;
        pixel_data[37][87] = 0;
        pixel_data[37][88] = 0;
        pixel_data[37][89] = 0;
        pixel_data[37][90] = 0;
        pixel_data[37][91] = 0;
        pixel_data[37][92] = 0;
        pixel_data[37][93] = 0;
        pixel_data[37][94] = 0;
        pixel_data[37][95] = 0;
        pixel_data[37][96] = 0;
        pixel_data[37][97] = 0;
        pixel_data[37][98] = 0;
        pixel_data[37][99] = 0; // y=37
        pixel_data[38][0] = 0;
        pixel_data[38][1] = 0;
        pixel_data[38][2] = 0;
        pixel_data[38][3] = 0;
        pixel_data[38][4] = 0;
        pixel_data[38][5] = 0;
        pixel_data[38][6] = 0;
        pixel_data[38][7] = 0;
        pixel_data[38][8] = 0;
        pixel_data[38][9] = 0;
        pixel_data[38][10] = 0;
        pixel_data[38][11] = 0;
        pixel_data[38][12] = 0;
        pixel_data[38][13] = 15;
        pixel_data[38][14] = 7;
        pixel_data[38][15] = 8;
        pixel_data[38][16] = 6;
        pixel_data[38][17] = 6;
        pixel_data[38][18] = 6;
        pixel_data[38][19] = 8;
        pixel_data[38][20] = 8;
        pixel_data[38][21] = 9;
        pixel_data[38][22] = 9;
        pixel_data[38][23] = 9;
        pixel_data[38][24] = 10;
        pixel_data[38][25] = 10;
        pixel_data[38][26] = 10;
        pixel_data[38][27] = 11;
        pixel_data[38][28] = 11;
        pixel_data[38][29] = 10;
        pixel_data[38][30] = 10;
        pixel_data[38][31] = 10;
        pixel_data[38][32] = 10;
        pixel_data[38][33] = 10;
        pixel_data[38][34] = 10;
        pixel_data[38][35] = 10;
        pixel_data[38][36] = 9;
        pixel_data[38][37] = 9;
        pixel_data[38][38] = 9;
        pixel_data[38][39] = 8;
        pixel_data[38][40] = 6;
        pixel_data[38][41] = 4;
        pixel_data[38][42] = 4;
        pixel_data[38][43] = 4;
        pixel_data[38][44] = 4;
        pixel_data[38][45] = 3;
        pixel_data[38][46] = 3;
        pixel_data[38][47] = 3;
        pixel_data[38][48] = 3;
        pixel_data[38][49] = 3;
        pixel_data[38][50] = 3;
        pixel_data[38][51] = 3;
        pixel_data[38][52] = 3;
        pixel_data[38][53] = 3;
        pixel_data[38][54] = 3;
        pixel_data[38][55] = 3;
        pixel_data[38][56] = 3;
        pixel_data[38][57] = 4;
        pixel_data[38][58] = 4;
        pixel_data[38][59] = 3;
        pixel_data[38][60] = 3;
        pixel_data[38][61] = 3;
        pixel_data[38][62] = 5;
        pixel_data[38][63] = 3;
        pixel_data[38][64] = 5;
        pixel_data[38][65] = 15;
        pixel_data[38][66] = 2;
        pixel_data[38][67] = 7;
        pixel_data[38][68] = 15;
        pixel_data[38][69] = 1;
        pixel_data[38][70] = 13;
        pixel_data[38][71] = 0;
        pixel_data[38][72] = 0;
        pixel_data[38][73] = 0;
        pixel_data[38][74] = 0;
        pixel_data[38][75] = 0;
        pixel_data[38][76] = 0;
        pixel_data[38][77] = 0;
        pixel_data[38][78] = 1;
        pixel_data[38][79] = 1;
        pixel_data[38][80] = 1;
        pixel_data[38][81] = 1;
        pixel_data[38][82] = 1;
        pixel_data[38][83] = 1;
        pixel_data[38][84] = 1;
        pixel_data[38][85] = 13;
        pixel_data[38][86] = 0;
        pixel_data[38][87] = 0;
        pixel_data[38][88] = 0;
        pixel_data[38][89] = 0;
        pixel_data[38][90] = 0;
        pixel_data[38][91] = 0;
        pixel_data[38][92] = 0;
        pixel_data[38][93] = 0;
        pixel_data[38][94] = 0;
        pixel_data[38][95] = 0;
        pixel_data[38][96] = 0;
        pixel_data[38][97] = 0;
        pixel_data[38][98] = 0;
        pixel_data[38][99] = 0; // y=38
        pixel_data[39][0] = 0;
        pixel_data[39][1] = 0;
        pixel_data[39][2] = 0;
        pixel_data[39][3] = 0;
        pixel_data[39][4] = 0;
        pixel_data[39][5] = 0;
        pixel_data[39][6] = 0;
        pixel_data[39][7] = 0;
        pixel_data[39][8] = 0;
        pixel_data[39][9] = 0;
        pixel_data[39][10] = 0;
        pixel_data[39][11] = 0;
        pixel_data[39][12] = 0;
        pixel_data[39][13] = 0;
        pixel_data[39][14] = 0;
        pixel_data[39][15] = 0;
        pixel_data[39][16] = 14;
        pixel_data[39][17] = 7;
        pixel_data[39][18] = 8;
        pixel_data[39][19] = 8;
        pixel_data[39][20] = 9;
        pixel_data[39][21] = 9;
        pixel_data[39][22] = 9;
        pixel_data[39][23] = 9;
        pixel_data[39][24] = 9;
        pixel_data[39][25] = 10;
        pixel_data[39][26] = 10;
        pixel_data[39][27] = 11;
        pixel_data[39][28] = 11;
        pixel_data[39][29] = 11;
        pixel_data[39][30] = 10;
        pixel_data[39][31] = 10;
        pixel_data[39][32] = 10;
        pixel_data[39][33] = 10;
        pixel_data[39][34] = 10;
        pixel_data[39][35] = 10;
        pixel_data[39][36] = 10;
        pixel_data[39][37] = 9;
        pixel_data[39][38] = 9;
        pixel_data[39][39] = 9;
        pixel_data[39][40] = 8;
        pixel_data[39][41] = 6;
        pixel_data[39][42] = 6;
        pixel_data[39][43] = 4;
        pixel_data[39][44] = 4;
        pixel_data[39][45] = 4;
        pixel_data[39][46] = 4;
        pixel_data[39][47] = 4;
        pixel_data[39][48] = 3;
        pixel_data[39][49] = 3;
        pixel_data[39][50] = 3;
        pixel_data[39][51] = 3;
        pixel_data[39][52] = 3;
        pixel_data[39][53] = 3;
        pixel_data[39][54] = 3;
        pixel_data[39][55] = 3;
        pixel_data[39][56] = 3;
        pixel_data[39][57] = 3;
        pixel_data[39][58] = 3;
        pixel_data[39][59] = 3;
        pixel_data[39][60] = 3;
        pixel_data[39][61] = 3;
        pixel_data[39][62] = 3;
        pixel_data[39][63] = 3;
        pixel_data[39][64] = 3;
        pixel_data[39][65] = 3;
        pixel_data[39][66] = 3;
        pixel_data[39][67] = 4;
        pixel_data[39][68] = 4;
        pixel_data[39][69] = 10;
        pixel_data[39][70] = 7;
        pixel_data[39][71] = 10;
        pixel_data[39][72] = 12;
        pixel_data[39][73] = 7;
        pixel_data[39][74] = 12;
        pixel_data[39][75] = 5;
        pixel_data[39][76] = 5;
        pixel_data[39][77] = 7;
        pixel_data[39][78] = 7;
        pixel_data[39][79] = 7;
        pixel_data[39][80] = 7;
        pixel_data[39][81] = 3;
        pixel_data[39][82] = 2;
        pixel_data[39][83] = 2;
        pixel_data[39][84] = 2;
        pixel_data[39][85] = 5;
        pixel_data[39][86] = 7;
        pixel_data[39][87] = 7;
        pixel_data[39][88] = 11;
        pixel_data[39][89] = 5;
        pixel_data[39][90] = 7;
        pixel_data[39][91] = 15;
        pixel_data[39][92] = 0;
        pixel_data[39][93] = 0;
        pixel_data[39][94] = 0;
        pixel_data[39][95] = 0;
        pixel_data[39][96] = 0;
        pixel_data[39][97] = 0;
        pixel_data[39][98] = 0;
        pixel_data[39][99] = 0; // y=39
        pixel_data[40][0] = 0;
        pixel_data[40][1] = 0;
        pixel_data[40][2] = 0;
        pixel_data[40][3] = 0;
        pixel_data[40][4] = 0;
        pixel_data[40][5] = 0;
        pixel_data[40][6] = 0;
        pixel_data[40][7] = 0;
        pixel_data[40][8] = 0;
        pixel_data[40][9] = 0;
        pixel_data[40][10] = 0;
        pixel_data[40][11] = 0;
        pixel_data[40][12] = 0;
        pixel_data[40][13] = 0;
        pixel_data[40][14] = 0;
        pixel_data[40][15] = 0;
        pixel_data[40][16] = 0;
        pixel_data[40][17] = 1;
        pixel_data[40][18] = 11;
        pixel_data[40][19] = 8;
        pixel_data[40][20] = 10;
        pixel_data[40][21] = 10;
        pixel_data[40][22] = 9;
        pixel_data[40][23] = 9;
        pixel_data[40][24] = 9;
        pixel_data[40][25] = 9;
        pixel_data[40][26] = 9;
        pixel_data[40][27] = 10;
        pixel_data[40][28] = 11;
        pixel_data[40][29] = 11;
        pixel_data[40][30] = 11;
        pixel_data[40][31] = 10;
        pixel_data[40][32] = 10;
        pixel_data[40][33] = 10;
        pixel_data[40][34] = 10;
        pixel_data[40][35] = 10;
        pixel_data[40][36] = 10;
        pixel_data[40][37] = 10;
        pixel_data[40][38] = 9;
        pixel_data[40][39] = 9;
        pixel_data[40][40] = 9;
        pixel_data[40][41] = 9;
        pixel_data[40][42] = 9;
        pixel_data[40][43] = 8;
        pixel_data[40][44] = 8;
        pixel_data[40][45] = 6;
        pixel_data[40][46] = 6;
        pixel_data[40][47] = 6;
        pixel_data[40][48] = 4;
        pixel_data[40][49] = 4;
        pixel_data[40][50] = 4;
        pixel_data[40][51] = 4;
        pixel_data[40][52] = 4;
        pixel_data[40][53] = 4;
        pixel_data[40][54] = 4;
        pixel_data[40][55] = 4;
        pixel_data[40][56] = 4;
        pixel_data[40][57] = 3;
        pixel_data[40][58] = 3;
        pixel_data[40][59] = 3;
        pixel_data[40][60] = 3;
        pixel_data[40][61] = 3;
        pixel_data[40][62] = 3;
        pixel_data[40][63] = 3;
        pixel_data[40][64] = 3;
        pixel_data[40][65] = 3;
        pixel_data[40][66] = 3;
        pixel_data[40][67] = 3;
        pixel_data[40][68] = 3;
        pixel_data[40][69] = 3;
        pixel_data[40][70] = 4;
        pixel_data[40][71] = 4;
        pixel_data[40][72] = 9;
        pixel_data[40][73] = 10;
        pixel_data[40][74] = 9;
        pixel_data[40][75] = 9;
        pixel_data[40][76] = 9;
        pixel_data[40][77] = 8;
        pixel_data[40][78] = 5;
        pixel_data[40][79] = 6;
        pixel_data[40][80] = 4;
        pixel_data[40][81] = 5;
        pixel_data[40][82] = 6;
        pixel_data[40][83] = 6;
        pixel_data[40][84] = 6;
        pixel_data[40][85] = 8;
        pixel_data[40][86] = 8;
        pixel_data[40][87] = 8;
        pixel_data[40][88] = 8;
        pixel_data[40][89] = 9;
        pixel_data[40][90] = 4;
        pixel_data[40][91] = 10;
        pixel_data[40][92] = 7;
        pixel_data[40][93] = 12;
        pixel_data[40][94] = 0;
        pixel_data[40][95] = 0;
        pixel_data[40][96] = 0;
        pixel_data[40][97] = 0;
        pixel_data[40][98] = 0;
        pixel_data[40][99] = 0; // y=40
        pixel_data[41][0] = 0;
        pixel_data[41][1] = 0;
        pixel_data[41][2] = 0;
        pixel_data[41][3] = 0;
        pixel_data[41][4] = 0;
        pixel_data[41][5] = 0;
        pixel_data[41][6] = 0;
        pixel_data[41][7] = 0;
        pixel_data[41][8] = 0;
        pixel_data[41][9] = 0;
        pixel_data[41][10] = 0;
        pixel_data[41][11] = 0;
        pixel_data[41][12] = 0;
        pixel_data[41][13] = 0;
        pixel_data[41][14] = 0;
        pixel_data[41][15] = 0;
        pixel_data[41][16] = 0;
        pixel_data[41][17] = 0;
        pixel_data[41][18] = 1;
        pixel_data[41][19] = 12;
        pixel_data[41][20] = 7;
        pixel_data[41][21] = 8;
        pixel_data[41][22] = 10;
        pixel_data[41][23] = 10;
        pixel_data[41][24] = 9;
        pixel_data[41][25] = 9;
        pixel_data[41][26] = 9;
        pixel_data[41][27] = 10;
        pixel_data[41][28] = 10;
        pixel_data[41][29] = 11;
        pixel_data[41][30] = 11;
        pixel_data[41][31] = 11;
        pixel_data[41][32] = 10;
        pixel_data[41][33] = 10;
        pixel_data[41][34] = 10;
        pixel_data[41][35] = 10;
        pixel_data[41][36] = 10;
        pixel_data[41][37] = 10;
        pixel_data[41][38] = 10;
        pixel_data[41][39] = 10;
        pixel_data[41][40] = 10;
        pixel_data[41][41] = 10;
        pixel_data[41][42] = 10;
        pixel_data[41][43] = 10;
        pixel_data[41][44] = 9;
        pixel_data[41][45] = 9;
        pixel_data[41][46] = 9;
        pixel_data[41][47] = 9;
        pixel_data[41][48] = 9;
        pixel_data[41][49] = 8;
        pixel_data[41][50] = 8;
        pixel_data[41][51] = 6;
        pixel_data[41][52] = 6;
        pixel_data[41][53] = 6;
        pixel_data[41][54] = 6;
        pixel_data[41][55] = 6;
        pixel_data[41][56] = 4;
        pixel_data[41][57] = 4;
        pixel_data[41][58] = 4;
        pixel_data[41][59] = 4;
        pixel_data[41][60] = 4;
        pixel_data[41][61] = 4;
        pixel_data[41][62] = 3;
        pixel_data[41][63] = 3;
        pixel_data[41][64] = 3;
        pixel_data[41][65] = 3;
        pixel_data[41][66] = 3;
        pixel_data[41][67] = 3;
        pixel_data[41][68] = 3;
        pixel_data[41][69] = 3;
        pixel_data[41][70] = 3;
        pixel_data[41][71] = 3;
        pixel_data[41][72] = 3;
        pixel_data[41][73] = 4;
        pixel_data[41][74] = 6;
        pixel_data[41][75] = 6;
        pixel_data[41][76] = 8;
        pixel_data[41][77] = 8;
        pixel_data[41][78] = 9;
        pixel_data[41][79] = 9;
        pixel_data[41][80] = 9;
        pixel_data[41][81] = 10;
        pixel_data[41][82] = 9;
        pixel_data[41][83] = 10;
        pixel_data[41][84] = 10;
        pixel_data[41][85] = 10;
        pixel_data[41][86] = 10;
        pixel_data[41][87] = 10;
        pixel_data[41][88] = 10;
        pixel_data[41][89] = 9;
        pixel_data[41][90] = 9;
        pixel_data[41][91] = 8;
        pixel_data[41][92] = 6;
        pixel_data[41][93] = 5;
        pixel_data[41][94] = 5;
        pixel_data[41][95] = 0;
        pixel_data[41][96] = 0;
        pixel_data[41][97] = 0;
        pixel_data[41][98] = 0;
        pixel_data[41][99] = 0; // y=41
        pixel_data[42][0] = 0;
        pixel_data[42][1] = 0;
        pixel_data[42][2] = 0;
        pixel_data[42][3] = 0;
        pixel_data[42][4] = 0;
        pixel_data[42][5] = 0;
        pixel_data[42][6] = 0;
        pixel_data[42][7] = 0;
        pixel_data[42][8] = 0;
        pixel_data[42][9] = 0;
        pixel_data[42][10] = 0;
        pixel_data[42][11] = 0;
        pixel_data[42][12] = 0;
        pixel_data[42][13] = 0;
        pixel_data[42][14] = 0;
        pixel_data[42][15] = 0;
        pixel_data[42][16] = 0;
        pixel_data[42][17] = 0;
        pixel_data[42][18] = 0;
        pixel_data[42][19] = 0;
        pixel_data[42][20] = 1;
        pixel_data[42][21] = 2;
        pixel_data[42][22] = 7;
        pixel_data[42][23] = 9;
        pixel_data[42][24] = 8;
        pixel_data[42][25] = 9;
        pixel_data[42][26] = 9;
        pixel_data[42][27] = 10;
        pixel_data[42][28] = 10;
        pixel_data[42][29] = 11;
        pixel_data[42][30] = 11;
        pixel_data[42][31] = 11;
        pixel_data[42][32] = 11;
        pixel_data[42][33] = 11;
        pixel_data[42][34] = 11;
        pixel_data[42][35] = 10;
        pixel_data[42][36] = 10;
        pixel_data[42][37] = 10;
        pixel_data[42][38] = 10;
        pixel_data[42][39] = 11;
        pixel_data[42][40] = 11;
        pixel_data[42][41] = 11;
        pixel_data[42][42] = 11;
        pixel_data[42][43] = 11;
        pixel_data[42][44] = 11;
        pixel_data[42][45] = 11;
        pixel_data[42][46] = 10;
        pixel_data[42][47] = 10;
        pixel_data[42][48] = 10;
        pixel_data[42][49] = 10;
        pixel_data[42][50] = 10;
        pixel_data[42][51] = 10;
        pixel_data[42][52] = 9;
        pixel_data[42][53] = 9;
        pixel_data[42][54] = 9;
        pixel_data[42][55] = 9;
        pixel_data[42][56] = 9;
        pixel_data[42][57] = 8;
        pixel_data[42][58] = 6;
        pixel_data[42][59] = 6;
        pixel_data[42][60] = 6;
        pixel_data[42][61] = 4;
        pixel_data[42][62] = 4;
        pixel_data[42][63] = 4;
        pixel_data[42][64] = 4;
        pixel_data[42][65] = 4;
        pixel_data[42][66] = 4;
        pixel_data[42][67] = 4;
        pixel_data[42][68] = 4;
        pixel_data[42][69] = 4;
        pixel_data[42][70] = 4;
        pixel_data[42][71] = 4;
        pixel_data[42][72] = 4;
        pixel_data[42][73] = 4;
        pixel_data[42][74] = 4;
        pixel_data[42][75] = 4;
        pixel_data[42][76] = 4;
        pixel_data[42][77] = 4;
        pixel_data[42][78] = 6;
        pixel_data[42][79] = 8;
        pixel_data[42][80] = 8;
        pixel_data[42][81] = 9;
        pixel_data[42][82] = 9;
        pixel_data[42][83] = 9;
        pixel_data[42][84] = 9;
        pixel_data[42][85] = 9;
        pixel_data[42][86] = 9;
        pixel_data[42][87] = 10;
        pixel_data[42][88] = 10;
        pixel_data[42][89] = 10;
        pixel_data[42][90] = 10;
        pixel_data[42][91] = 10;
        pixel_data[42][92] = 9;
        pixel_data[42][93] = 8;
        pixel_data[42][94] = 8;
        pixel_data[42][95] = 7;
        pixel_data[42][96] = 12;
        pixel_data[42][97] = 12;
        pixel_data[42][98] = 7;
        pixel_data[42][99] = 1; // y=42
        pixel_data[43][0] = 0;
        pixel_data[43][1] = 0;
        pixel_data[43][2] = 0;
        pixel_data[43][3] = 0;
        pixel_data[43][4] = 0;
        pixel_data[43][5] = 0;
        pixel_data[43][6] = 0;
        pixel_data[43][7] = 0;
        pixel_data[43][8] = 0;
        pixel_data[43][9] = 0;
        pixel_data[43][10] = 0;
        pixel_data[43][11] = 0;
        pixel_data[43][12] = 0;
        pixel_data[43][13] = 0;
        pixel_data[43][14] = 0;
        pixel_data[43][15] = 0;
        pixel_data[43][16] = 0;
        pixel_data[43][17] = 0;
        pixel_data[43][18] = 0;
        pixel_data[43][19] = 15;
        pixel_data[43][20] = 10;
        pixel_data[43][21] = 8;
        pixel_data[43][22] = 8;
        pixel_data[43][23] = 8;
        pixel_data[43][24] = 9;
        pixel_data[43][25] = 10;
        pixel_data[43][26] = 10;
        pixel_data[43][27] = 11;
        pixel_data[43][28] = 11;
        pixel_data[43][29] = 11;
        pixel_data[43][30] = 11;
        pixel_data[43][31] = 11;
        pixel_data[43][32] = 11;
        pixel_data[43][33] = 11;
        pixel_data[43][34] = 11;
        pixel_data[43][35] = 11;
        pixel_data[43][36] = 11;
        pixel_data[43][37] = 11;
        pixel_data[43][38] = 11;
        pixel_data[43][39] = 11;
        pixel_data[43][40] = 12;
        pixel_data[43][41] = 12;
        pixel_data[43][42] = 11;
        pixel_data[43][43] = 11;
        pixel_data[43][44] = 11;
        pixel_data[43][45] = 11;
        pixel_data[43][46] = 11;
        pixel_data[43][47] = 11;
        pixel_data[43][48] = 11;
        pixel_data[43][49] = 11;
        pixel_data[43][50] = 11;
        pixel_data[43][51] = 10;
        pixel_data[43][52] = 10;
        pixel_data[43][53] = 10;
        pixel_data[43][54] = 10;
        pixel_data[43][55] = 10;
        pixel_data[43][56] = 10;
        pixel_data[43][57] = 10;
        pixel_data[43][58] = 9;
        pixel_data[43][59] = 9;
        pixel_data[43][60] = 9;
        pixel_data[43][61] = 8;
        pixel_data[43][62] = 8;
        pixel_data[43][63] = 8;
        pixel_data[43][64] = 8;
        pixel_data[43][65] = 6;
        pixel_data[43][66] = 6;
        pixel_data[43][67] = 6;
        pixel_data[43][68] = 6;
        pixel_data[43][69] = 6;
        pixel_data[43][70] = 6;
        pixel_data[43][71] = 6;
        pixel_data[43][72] = 6;
        pixel_data[43][73] = 6;
        pixel_data[43][74] = 6;
        pixel_data[43][75] = 6;
        pixel_data[43][76] = 6;
        pixel_data[43][77] = 6;
        pixel_data[43][78] = 6;
        pixel_data[43][79] = 6;
        pixel_data[43][80] = 6;
        pixel_data[43][81] = 4;
        pixel_data[43][82] = 6;
        pixel_data[43][83] = 6;
        pixel_data[43][84] = 8;
        pixel_data[43][85] = 8;
        pixel_data[43][86] = 8;
        pixel_data[43][87] = 9;
        pixel_data[43][88] = 9;
        pixel_data[43][89] = 10;
        pixel_data[43][90] = 10;
        pixel_data[43][91] = 11;
        pixel_data[43][92] = 10;
        pixel_data[43][93] = 9;
        pixel_data[43][94] = 8;
        pixel_data[43][95] = 9;
        pixel_data[43][96] = 11;
        pixel_data[43][97] = 11;
        pixel_data[43][98] = 11;
        pixel_data[43][99] = 7; // y=43
        pixel_data[44][0] = 0;
        pixel_data[44][1] = 0;
        pixel_data[44][2] = 0;
        pixel_data[44][3] = 0;
        pixel_data[44][4] = 0;
        pixel_data[44][5] = 0;
        pixel_data[44][6] = 0;
        pixel_data[44][7] = 0;
        pixel_data[44][8] = 0;
        pixel_data[44][9] = 0;
        pixel_data[44][10] = 0;
        pixel_data[44][11] = 0;
        pixel_data[44][12] = 0;
        pixel_data[44][13] = 0;
        pixel_data[44][14] = 0;
        pixel_data[44][15] = 0;
        pixel_data[44][16] = 0;
        pixel_data[44][17] = 15;
        pixel_data[44][18] = 5;
        pixel_data[44][19] = 6;
        pixel_data[44][20] = 8;
        pixel_data[44][21] = 8;
        pixel_data[44][22] = 8;
        pixel_data[44][23] = 9;
        pixel_data[44][24] = 10;
        pixel_data[44][25] = 11;
        pixel_data[44][26] = 11;
        pixel_data[44][27] = 11;
        pixel_data[44][28] = 11;
        pixel_data[44][29] = 12;
        pixel_data[44][30] = 12;
        pixel_data[44][31] = 12;
        pixel_data[44][32] = 12;
        pixel_data[44][33] = 12;
        pixel_data[44][34] = 12;
        pixel_data[44][35] = 11;
        pixel_data[44][36] = 11;
        pixel_data[44][37] = 11;
        pixel_data[44][38] = 12;
        pixel_data[44][39] = 12;
        pixel_data[44][40] = 12;
        pixel_data[44][41] = 12;
        pixel_data[44][42] = 12;
        pixel_data[44][43] = 12;
        pixel_data[44][44] = 12;
        pixel_data[44][45] = 12;
        pixel_data[44][46] = 11;
        pixel_data[44][47] = 11;
        pixel_data[44][48] = 11;
        pixel_data[44][49] = 11;
        pixel_data[44][50] = 11;
        pixel_data[44][51] = 11;
        pixel_data[44][52] = 11;
        pixel_data[44][53] = 11;
        pixel_data[44][54] = 11;
        pixel_data[44][55] = 11;
        pixel_data[44][56] = 10;
        pixel_data[44][57] = 10;
        pixel_data[44][58] = 10;
        pixel_data[44][59] = 10;
        pixel_data[44][60] = 10;
        pixel_data[44][61] = 10;
        pixel_data[44][62] = 9;
        pixel_data[44][63] = 9;
        pixel_data[44][64] = 9;
        pixel_data[44][65] = 9;
        pixel_data[44][66] = 9;
        pixel_data[44][67] = 9;
        pixel_data[44][68] = 9;
        pixel_data[44][69] = 9;
        pixel_data[44][70] = 9;
        pixel_data[44][71] = 9;
        pixel_data[44][72] = 9;
        pixel_data[44][73] = 8;
        pixel_data[44][74] = 9;
        pixel_data[44][75] = 9;
        pixel_data[44][76] = 8;
        pixel_data[44][77] = 8;
        pixel_data[44][78] = 8;
        pixel_data[44][79] = 6;
        pixel_data[44][80] = 6;
        pixel_data[44][81] = 6;
        pixel_data[44][82] = 6;
        pixel_data[44][83] = 6;
        pixel_data[44][84] = 6;
        pixel_data[44][85] = 8;
        pixel_data[44][86] = 8;
        pixel_data[44][87] = 8;
        pixel_data[44][88] = 9;
        pixel_data[44][89] = 9;
        pixel_data[44][90] = 10;
        pixel_data[44][91] = 11;
        pixel_data[44][92] = 11;
        pixel_data[44][93] = 10;
        pixel_data[44][94] = 9;
        pixel_data[44][95] = 9;
        pixel_data[44][96] = 10;
        pixel_data[44][97] = 11;
        pixel_data[44][98] = 11;
        pixel_data[44][99] = 11; // y=44
        pixel_data[45][0] = 0;
        pixel_data[45][1] = 0;
        pixel_data[45][2] = 0;
        pixel_data[45][3] = 0;
        pixel_data[45][4] = 0;
        pixel_data[45][5] = 0;
        pixel_data[45][6] = 0;
        pixel_data[45][7] = 0;
        pixel_data[45][8] = 0;
        pixel_data[45][9] = 0;
        pixel_data[45][10] = 0;
        pixel_data[45][11] = 0;
        pixel_data[45][12] = 0;
        pixel_data[45][13] = 0;
        pixel_data[45][14] = 0;
        pixel_data[45][15] = 1;
        pixel_data[45][16] = 11;
        pixel_data[45][17] = 8;
        pixel_data[45][18] = 8;
        pixel_data[45][19] = 6;
        pixel_data[45][20] = 8;
        pixel_data[45][21] = 9;
        pixel_data[45][22] = 10;
        pixel_data[45][23] = 11;
        pixel_data[45][24] = 11;
        pixel_data[45][25] = 12;
        pixel_data[45][26] = 12;
        pixel_data[45][27] = 12;
        pixel_data[45][28] = 12;
        pixel_data[45][29] = 12;
        pixel_data[45][30] = 12;
        pixel_data[45][31] = 12;
        pixel_data[45][32] = 13;
        pixel_data[45][33] = 13;
        pixel_data[45][34] = 12;
        pixel_data[45][35] = 12;
        pixel_data[45][36] = 11;
        pixel_data[45][37] = 12;
        pixel_data[45][38] = 12;
        pixel_data[45][39] = 12;
        pixel_data[45][40] = 12;
        pixel_data[45][41] = 12;
        pixel_data[45][42] = 12;
        pixel_data[45][43] = 12;
        pixel_data[45][44] = 12;
        pixel_data[45][45] = 12;
        pixel_data[45][46] = 12;
        pixel_data[45][47] = 12;
        pixel_data[45][48] = 12;
        pixel_data[45][49] = 12;
        pixel_data[45][50] = 12;
        pixel_data[45][51] = 11;
        pixel_data[45][52] = 11;
        pixel_data[45][53] = 11;
        pixel_data[45][54] = 11;
        pixel_data[45][55] = 11;
        pixel_data[45][56] = 11;
        pixel_data[45][57] = 11;
        pixel_data[45][58] = 10;
        pixel_data[45][59] = 10;
        pixel_data[45][60] = 10;
        pixel_data[45][61] = 10;
        pixel_data[45][62] = 10;
        pixel_data[45][63] = 10;
        pixel_data[45][64] = 10;
        pixel_data[45][65] = 10;
        pixel_data[45][66] = 9;
        pixel_data[45][67] = 9;
        pixel_data[45][68] = 9;
        pixel_data[45][69] = 9;
        pixel_data[45][70] = 9;
        pixel_data[45][71] = 9;
        pixel_data[45][72] = 9;
        pixel_data[45][73] = 9;
        pixel_data[45][74] = 9;
        pixel_data[45][75] = 9;
        pixel_data[45][76] = 9;
        pixel_data[45][77] = 9;
        pixel_data[45][78] = 9;
        pixel_data[45][79] = 8;
        pixel_data[45][80] = 8;
        pixel_data[45][81] = 8;
        pixel_data[45][82] = 6;
        pixel_data[45][83] = 6;
        pixel_data[45][84] = 6;
        pixel_data[45][85] = 6;
        pixel_data[45][86] = 8;
        pixel_data[45][87] = 8;
        pixel_data[45][88] = 9;
        pixel_data[45][89] = 9;
        pixel_data[45][90] = 10;
        pixel_data[45][91] = 11;
        pixel_data[45][92] = 11;
        pixel_data[45][93] = 10;
        pixel_data[45][94] = 10;
        pixel_data[45][95] = 9;
        pixel_data[45][96] = 10;
        pixel_data[45][97] = 11;
        pixel_data[45][98] = 11;
        pixel_data[45][99] = 11; // y=45
        pixel_data[46][0] = 0;
        pixel_data[46][1] = 0;
        pixel_data[46][2] = 0;
        pixel_data[46][3] = 0;
        pixel_data[46][4] = 0;
        pixel_data[46][5] = 0;
        pixel_data[46][6] = 0;
        pixel_data[46][7] = 0;
        pixel_data[46][8] = 0;
        pixel_data[46][9] = 0;
        pixel_data[46][10] = 0;
        pixel_data[46][11] = 0;
        pixel_data[46][12] = 0;
        pixel_data[46][13] = 1;
        pixel_data[46][14] = 7;
        pixel_data[46][15] = 6;
        pixel_data[46][16] = 8;
        pixel_data[46][17] = 6;
        pixel_data[46][18] = 8;
        pixel_data[46][19] = 9;
        pixel_data[46][20] = 10;
        pixel_data[46][21] = 11;
        pixel_data[46][22] = 11;
        pixel_data[46][23] = 12;
        pixel_data[46][24] = 12;
        pixel_data[46][25] = 12;
        pixel_data[46][26] = 12;
        pixel_data[46][27] = 12;
        pixel_data[46][28] = 12;
        pixel_data[46][29] = 12;
        pixel_data[46][30] = 12;
        pixel_data[46][31] = 13;
        pixel_data[46][32] = 13;
        pixel_data[46][33] = 13;
        pixel_data[46][34] = 12;
        pixel_data[46][35] = 12;
        pixel_data[46][36] = 12;
        pixel_data[46][37] = 12;
        pixel_data[46][38] = 12;
        pixel_data[46][39] = 12;
        pixel_data[46][40] = 12;
        pixel_data[46][41] = 13;
        pixel_data[46][42] = 12;
        pixel_data[46][43] = 12;
        pixel_data[46][44] = 12;
        pixel_data[46][45] = 12;
        pixel_data[46][46] = 12;
        pixel_data[46][47] = 12;
        pixel_data[46][48] = 12;
        pixel_data[46][49] = 12;
        pixel_data[46][50] = 12;
        pixel_data[46][51] = 12;
        pixel_data[46][52] = 12;
        pixel_data[46][53] = 11;
        pixel_data[46][54] = 11;
        pixel_data[46][55] = 11;
        pixel_data[46][56] = 11;
        pixel_data[46][57] = 11;
        pixel_data[46][58] = 11;
        pixel_data[46][59] = 11;
        pixel_data[46][60] = 10;
        pixel_data[46][61] = 10;
        pixel_data[46][62] = 10;
        pixel_data[46][63] = 10;
        pixel_data[46][64] = 10;
        pixel_data[46][65] = 10;
        pixel_data[46][66] = 10;
        pixel_data[46][67] = 10;
        pixel_data[46][68] = 10;
        pixel_data[46][69] = 10;
        pixel_data[46][70] = 10;
        pixel_data[46][71] = 10;
        pixel_data[46][72] = 10;
        pixel_data[46][73] = 10;
        pixel_data[46][74] = 9;
        pixel_data[46][75] = 9;
        pixel_data[46][76] = 9;
        pixel_data[46][77] = 9;
        pixel_data[46][78] = 9;
        pixel_data[46][79] = 9;
        pixel_data[46][80] = 9;
        pixel_data[46][81] = 9;
        pixel_data[46][82] = 8;
        pixel_data[46][83] = 8;
        pixel_data[46][84] = 8;
        pixel_data[46][85] = 8;
        pixel_data[46][86] = 6;
        pixel_data[46][87] = 6;
        pixel_data[46][88] = 8;
        pixel_data[46][89] = 9;
        pixel_data[46][90] = 10;
        pixel_data[46][91] = 11;
        pixel_data[46][92] = 11;
        pixel_data[46][93] = 11;
        pixel_data[46][94] = 10;
        pixel_data[46][95] = 9;
        pixel_data[46][96] = 10;
        pixel_data[46][97] = 10;
        pixel_data[46][98] = 11;
        pixel_data[46][99] = 11; // y=46
        pixel_data[47][0] = 0;
        pixel_data[47][1] = 0;
        pixel_data[47][2] = 0;
        pixel_data[47][3] = 0;
        pixel_data[47][4] = 0;
        pixel_data[47][5] = 0;
        pixel_data[47][6] = 0;
        pixel_data[47][7] = 0;
        pixel_data[47][8] = 0;
        pixel_data[47][9] = 0;
        pixel_data[47][10] = 0;
        pixel_data[47][11] = 15;
        pixel_data[47][12] = 7;
        pixel_data[47][13] = 8;
        pixel_data[47][14] = 8;
        pixel_data[47][15] = 8;
        pixel_data[47][16] = 8;
        pixel_data[47][17] = 9;
        pixel_data[47][18] = 10;
        pixel_data[47][19] = 11;
        pixel_data[47][20] = 12;
        pixel_data[47][21] = 12;
        pixel_data[47][22] = 12;
        pixel_data[47][23] = 12;
        pixel_data[47][24] = 12;
        pixel_data[47][25] = 12;
        pixel_data[47][26] = 12;
        pixel_data[47][27] = 12;
        pixel_data[47][28] = 12;
        pixel_data[47][29] = 12;
        pixel_data[47][30] = 12;
        pixel_data[47][31] = 13;
        pixel_data[47][32] = 13;
        pixel_data[47][33] = 13;
        pixel_data[47][34] = 12;
        pixel_data[47][35] = 12;
        pixel_data[47][36] = 12;
        pixel_data[47][37] = 12;
        pixel_data[47][38] = 13;
        pixel_data[47][39] = 13;
        pixel_data[47][40] = 13;
        pixel_data[47][41] = 13;
        pixel_data[47][42] = 13;
        pixel_data[47][43] = 13;
        pixel_data[47][44] = 13;
        pixel_data[47][45] = 13;
        pixel_data[47][46] = 13;
        pixel_data[47][47] = 13;
        pixel_data[47][48] = 12;
        pixel_data[47][49] = 12;
        pixel_data[47][50] = 12;
        pixel_data[47][51] = 12;
        pixel_data[47][52] = 12;
        pixel_data[47][53] = 12;
        pixel_data[47][54] = 11;
        pixel_data[47][55] = 11;
        pixel_data[47][56] = 11;
        pixel_data[47][57] = 11;
        pixel_data[47][58] = 11;
        pixel_data[47][59] = 11;
        pixel_data[47][60] = 11;
        pixel_data[47][61] = 11;
        pixel_data[47][62] = 11;
        pixel_data[47][63] = 10;
        pixel_data[47][64] = 10;
        pixel_data[47][65] = 10;
        pixel_data[47][66] = 10;
        pixel_data[47][67] = 10;
        pixel_data[47][68] = 10;
        pixel_data[47][69] = 10;
        pixel_data[47][70] = 10;
        pixel_data[47][71] = 10;
        pixel_data[47][72] = 10;
        pixel_data[47][73] = 10;
        pixel_data[47][74] = 10;
        pixel_data[47][75] = 10;
        pixel_data[47][76] = 10;
        pixel_data[47][77] = 10;
        pixel_data[47][78] = 10;
        pixel_data[47][79] = 9;
        pixel_data[47][80] = 9;
        pixel_data[47][81] = 9;
        pixel_data[47][82] = 9;
        pixel_data[47][83] = 8;
        pixel_data[47][84] = 8;
        pixel_data[47][85] = 8;
        pixel_data[47][86] = 8;
        pixel_data[47][87] = 6;
        pixel_data[47][88] = 8;
        pixel_data[47][89] = 9;
        pixel_data[47][90] = 10;
        pixel_data[47][91] = 11;
        pixel_data[47][92] = 11;
        pixel_data[47][93] = 11;
        pixel_data[47][94] = 10;
        pixel_data[47][95] = 10;
        pixel_data[47][96] = 10;
        pixel_data[47][97] = 11;
        pixel_data[47][98] = 11;
        pixel_data[47][99] = 11; // y=47
        pixel_data[48][0] = 0;
        pixel_data[48][1] = 0;
        pixel_data[48][2] = 0;
        pixel_data[48][3] = 0;
        pixel_data[48][4] = 0;
        pixel_data[48][5] = 0;
        pixel_data[48][6] = 0;
        pixel_data[48][7] = 0;
        pixel_data[48][8] = 0;
        pixel_data[48][9] = 1;
        pixel_data[48][10] = 7;
        pixel_data[48][11] = 6;
        pixel_data[48][12] = 8;
        pixel_data[48][13] = 8;
        pixel_data[48][14] = 8;
        pixel_data[48][15] = 9;
        pixel_data[48][16] = 10;
        pixel_data[48][17] = 11;
        pixel_data[48][18] = 11;
        pixel_data[48][19] = 12;
        pixel_data[48][20] = 12;
        pixel_data[48][21] = 12;
        pixel_data[48][22] = 12;
        pixel_data[48][23] = 12;
        pixel_data[48][24] = 12;
        pixel_data[48][25] = 12;
        pixel_data[48][26] = 12;
        pixel_data[48][27] = 12;
        pixel_data[48][28] = 12;
        pixel_data[48][29] = 13;
        pixel_data[48][30] = 13;
        pixel_data[48][31] = 13;
        pixel_data[48][32] = 13;
        pixel_data[48][33] = 13;
        pixel_data[48][34] = 12;
        pixel_data[48][35] = 13;
        pixel_data[48][36] = 13;
        pixel_data[48][37] = 13;
        pixel_data[48][38] = 13;
        pixel_data[48][39] = 13;
        pixel_data[48][40] = 13;
        pixel_data[48][41] = 13;
        pixel_data[48][42] = 13;
        pixel_data[48][43] = 13;
        pixel_data[48][44] = 13;
        pixel_data[48][45] = 13;
        pixel_data[48][46] = 13;
        pixel_data[48][47] = 13;
        pixel_data[48][48] = 12;
        pixel_data[48][49] = 12;
        pixel_data[48][50] = 12;
        pixel_data[48][51] = 12;
        pixel_data[48][52] = 12;
        pixel_data[48][53] = 12;
        pixel_data[48][54] = 12;
        pixel_data[48][55] = 11;
        pixel_data[48][56] = 11;
        pixel_data[48][57] = 11;
        pixel_data[48][58] = 11;
        pixel_data[48][59] = 11;
        pixel_data[48][60] = 11;
        pixel_data[48][61] = 11;
        pixel_data[48][62] = 11;
        pixel_data[48][63] = 11;
        pixel_data[48][64] = 10;
        pixel_data[48][65] = 10;
        pixel_data[48][66] = 10;
        pixel_data[48][67] = 10;
        pixel_data[48][68] = 10;
        pixel_data[48][69] = 10;
        pixel_data[48][70] = 10;
        pixel_data[48][71] = 10;
        pixel_data[48][72] = 10;
        pixel_data[48][73] = 10;
        pixel_data[48][74] = 10;
        pixel_data[48][75] = 10;
        pixel_data[48][76] = 10;
        pixel_data[48][77] = 10;
        pixel_data[48][78] = 10;
        pixel_data[48][79] = 10;
        pixel_data[48][80] = 9;
        pixel_data[48][81] = 9;
        pixel_data[48][82] = 9;
        pixel_data[48][83] = 8;
        pixel_data[48][84] = 8;
        pixel_data[48][85] = 8;
        pixel_data[48][86] = 8;
        pixel_data[48][87] = 8;
        pixel_data[48][88] = 9;
        pixel_data[48][89] = 10;
        pixel_data[48][90] = 11;
        pixel_data[48][91] = 11;
        pixel_data[48][92] = 11;
        pixel_data[48][93] = 10;
        pixel_data[48][94] = 9;
        pixel_data[48][95] = 9;
        pixel_data[48][96] = 10;
        pixel_data[48][97] = 11;
        pixel_data[48][98] = 11;
        pixel_data[48][99] = 11; // y=48
        pixel_data[49][0] = 0;
        pixel_data[49][1] = 0;
        pixel_data[49][2] = 0;
        pixel_data[49][3] = 0;
        pixel_data[49][4] = 0;
        pixel_data[49][5] = 0;
        pixel_data[49][6] = 0;
        pixel_data[49][7] = 0;
        pixel_data[49][8] = 7;
        pixel_data[49][9] = 8;
        pixel_data[49][10] = 6;
        pixel_data[49][11] = 8;
        pixel_data[49][12] = 8;
        pixel_data[49][13] = 9;
        pixel_data[49][14] = 10;
        pixel_data[49][15] = 11;
        pixel_data[49][16] = 12;
        pixel_data[49][17] = 12;
        pixel_data[49][18] = 12;
        pixel_data[49][19] = 12;
        pixel_data[49][20] = 12;
        pixel_data[49][21] = 12;
        pixel_data[49][22] = 12;
        pixel_data[49][23] = 12;
        pixel_data[49][24] = 12;
        pixel_data[49][25] = 12;
        pixel_data[49][26] = 12;
        pixel_data[49][27] = 12;
        pixel_data[49][28] = 13;
        pixel_data[49][29] = 13;
        pixel_data[49][30] = 13;
        pixel_data[49][31] = 13;
        pixel_data[49][32] = 13;
        pixel_data[49][33] = 13;
        pixel_data[49][34] = 13;
        pixel_data[49][35] = 13;
        pixel_data[49][36] = 13;
        pixel_data[49][37] = 13;
        pixel_data[49][38] = 13;
        pixel_data[49][39] = 13;
        pixel_data[49][40] = 13;
        pixel_data[49][41] = 13;
        pixel_data[49][42] = 13;
        pixel_data[49][43] = 13;
        pixel_data[49][44] = 13;
        pixel_data[49][45] = 13;
        pixel_data[49][46] = 13;
        pixel_data[49][47] = 13;
        pixel_data[49][48] = 13;
        pixel_data[49][49] = 12;
        pixel_data[49][50] = 12;
        pixel_data[49][51] = 12;
        pixel_data[49][52] = 12;
        pixel_data[49][53] = 12;
        pixel_data[49][54] = 12;
        pixel_data[49][55] = 12;
        pixel_data[49][56] = 11;
        pixel_data[49][57] = 11;
        pixel_data[49][58] = 11;
        pixel_data[49][59] = 11;
        pixel_data[49][60] = 11;
        pixel_data[49][61] = 11;
        pixel_data[49][62] = 11;
        pixel_data[49][63] = 11;
        pixel_data[49][64] = 11;
        pixel_data[49][65] = 11;
        pixel_data[49][66] = 10;
        pixel_data[49][67] = 10;
        pixel_data[49][68] = 10;
        pixel_data[49][69] = 10;
        pixel_data[49][70] = 10;
        pixel_data[49][71] = 10;
        pixel_data[49][72] = 10;
        pixel_data[49][73] = 10;
        pixel_data[49][74] = 10;
        pixel_data[49][75] = 10;
        pixel_data[49][76] = 10;
        pixel_data[49][77] = 10;
        pixel_data[49][78] = 10;
        pixel_data[49][79] = 10;
        pixel_data[49][80] = 10;
        pixel_data[49][81] = 9;
        pixel_data[49][82] = 9;
        pixel_data[49][83] = 8;
        pixel_data[49][84] = 8;
        pixel_data[49][85] = 8;
        pixel_data[49][86] = 6;
        pixel_data[49][87] = 8;
        pixel_data[49][88] = 9;
        pixel_data[49][89] = 10;
        pixel_data[49][90] = 11;
        pixel_data[49][91] = 11;
        pixel_data[49][92] = 10;
        pixel_data[49][93] = 9;
        pixel_data[49][94] = 9;
        pixel_data[49][95] = 9;
        pixel_data[49][96] = 10;
        pixel_data[49][97] = 11;
        pixel_data[49][98] = 11;
        pixel_data[49][99] = 11; // y=49
        pixel_data[50][0] = 0;
        pixel_data[50][1] = 0;
        pixel_data[50][2] = 0;
        pixel_data[50][3] = 0;
        pixel_data[50][4] = 0;
        pixel_data[50][5] = 0;
        pixel_data[50][6] = 0;
        pixel_data[50][7] = 7;
        pixel_data[50][8] = 4;
        pixel_data[50][9] = 6;
        pixel_data[50][10] = 6;
        pixel_data[50][11] = 8;
        pixel_data[50][12] = 10;
        pixel_data[50][13] = 11;
        pixel_data[50][14] = 11;
        pixel_data[50][15] = 11;
        pixel_data[50][16] = 11;
        pixel_data[50][17] = 12;
        pixel_data[50][18] = 12;
        pixel_data[50][19] = 12;
        pixel_data[50][20] = 12;
        pixel_data[50][21] = 12;
        pixel_data[50][22] = 12;
        pixel_data[50][23] = 12;
        pixel_data[50][24] = 12;
        pixel_data[50][25] = 12;
        pixel_data[50][26] = 12;
        pixel_data[50][27] = 12;
        pixel_data[50][28] = 13;
        pixel_data[50][29] = 13;
        pixel_data[50][30] = 13;
        pixel_data[50][31] = 13;
        pixel_data[50][32] = 13;
        pixel_data[50][33] = 13;
        pixel_data[50][34] = 1;
        pixel_data[50][35] = 1;
        pixel_data[50][36] = 1;
        pixel_data[50][37] = 13;
        pixel_data[50][38] = 13;
        pixel_data[50][39] = 13;
        pixel_data[50][40] = 13;
        pixel_data[50][41] = 13;
        pixel_data[50][42] = 13;
        pixel_data[50][43] = 13;
        pixel_data[50][44] = 13;
        pixel_data[50][45] = 13;
        pixel_data[50][46] = 13;
        pixel_data[50][47] = 13;
        pixel_data[50][48] = 13;
        pixel_data[50][49] = 13;
        pixel_data[50][50] = 13;
        pixel_data[50][51] = 12;
        pixel_data[50][52] = 12;
        pixel_data[50][53] = 12;
        pixel_data[50][54] = 12;
        pixel_data[50][55] = 12;
        pixel_data[50][56] = 12;
        pixel_data[50][57] = 12;
        pixel_data[50][58] = 11;
        pixel_data[50][59] = 11;
        pixel_data[50][60] = 11;
        pixel_data[50][61] = 11;
        pixel_data[50][62] = 11;
        pixel_data[50][63] = 11;
        pixel_data[50][64] = 11;
        pixel_data[50][65] = 11;
        pixel_data[50][66] = 11;
        pixel_data[50][67] = 11;
        pixel_data[50][68] = 10;
        pixel_data[50][69] = 10;
        pixel_data[50][70] = 10;
        pixel_data[50][71] = 10;
        pixel_data[50][72] = 10;
        pixel_data[50][73] = 10;
        pixel_data[50][74] = 10;
        pixel_data[50][75] = 10;
        pixel_data[50][76] = 10;
        pixel_data[50][77] = 10;
        pixel_data[50][78] = 10;
        pixel_data[50][79] = 10;
        pixel_data[50][80] = 10;
        pixel_data[50][81] = 9;
        pixel_data[50][82] = 9;
        pixel_data[50][83] = 8;
        pixel_data[50][84] = 8;
        pixel_data[50][85] = 6;
        pixel_data[50][86] = 6;
        pixel_data[50][87] = 8;
        pixel_data[50][88] = 10;
        pixel_data[50][89] = 10;
        pixel_data[50][90] = 10;
        pixel_data[50][91] = 9;
        pixel_data[50][92] = 8;
        pixel_data[50][93] = 8;
        pixel_data[50][94] = 8;
        pixel_data[50][95] = 9;
        pixel_data[50][96] = 9;
        pixel_data[50][97] = 10;
        pixel_data[50][98] = 10;
        pixel_data[50][99] = 11; // y=50
        pixel_data[51][0] = 0;
        pixel_data[51][1] = 0;
        pixel_data[51][2] = 0;
        pixel_data[51][3] = 0;
        pixel_data[51][4] = 0;
        pixel_data[51][5] = 0;
        pixel_data[51][6] = 8;
        pixel_data[51][7] = 6;
        pixel_data[51][8] = 6;
        pixel_data[51][9] = 6;
        pixel_data[51][10] = 8;
        pixel_data[51][11] = 10;
        pixel_data[51][12] = 11;
        pixel_data[51][13] = 11;
        pixel_data[51][14] = 11;
        pixel_data[51][15] = 11;
        pixel_data[51][16] = 11;
        pixel_data[51][17] = 12;
        pixel_data[51][18] = 12;
        pixel_data[51][19] = 12;
        pixel_data[51][20] = 12;
        pixel_data[51][21] = 12;
        pixel_data[51][22] = 12;
        pixel_data[51][23] = 12;
        pixel_data[51][24] = 12;
        pixel_data[51][25] = 12;
        pixel_data[51][26] = 12;
        pixel_data[51][27] = 13;
        pixel_data[51][28] = 13;
        pixel_data[51][29] = 13;
        pixel_data[51][30] = 13;
        pixel_data[51][31] = 1;
        pixel_data[51][32] = 1;
        pixel_data[51][33] = 1;
        pixel_data[51][34] = 1;
        pixel_data[51][35] = 1;
        pixel_data[51][36] = 1;
        pixel_data[51][37] = 13;
        pixel_data[51][38] = 13;
        pixel_data[51][39] = 13;
        pixel_data[51][40] = 13;
        pixel_data[51][41] = 13;
        pixel_data[51][42] = 13;
        pixel_data[51][43] = 13;
        pixel_data[51][44] = 13;
        pixel_data[51][45] = 13;
        pixel_data[51][46] = 13;
        pixel_data[51][47] = 13;
        pixel_data[51][48] = 13;
        pixel_data[51][49] = 13;
        pixel_data[51][50] = 13;
        pixel_data[51][51] = 13;
        pixel_data[51][52] = 12;
        pixel_data[51][53] = 12;
        pixel_data[51][54] = 12;
        pixel_data[51][55] = 12;
        pixel_data[51][56] = 12;
        pixel_data[51][57] = 12;
        pixel_data[51][58] = 12;
        pixel_data[51][59] = 12;
        pixel_data[51][60] = 12;
        pixel_data[51][61] = 11;
        pixel_data[51][62] = 11;
        pixel_data[51][63] = 11;
        pixel_data[51][64] = 11;
        pixel_data[51][65] = 11;
        pixel_data[51][66] = 11;
        pixel_data[51][67] = 11;
        pixel_data[51][68] = 11;
        pixel_data[51][69] = 10;
        pixel_data[51][70] = 10;
        pixel_data[51][71] = 10;
        pixel_data[51][72] = 10;
        pixel_data[51][73] = 10;
        pixel_data[51][74] = 10;
        pixel_data[51][75] = 10;
        pixel_data[51][76] = 10;
        pixel_data[51][77] = 10;
        pixel_data[51][78] = 10;
        pixel_data[51][79] = 10;
        pixel_data[51][80] = 9;
        pixel_data[51][81] = 9;
        pixel_data[51][82] = 8;
        pixel_data[51][83] = 8;
        pixel_data[51][84] = 6;
        pixel_data[51][85] = 6;
        pixel_data[51][86] = 8;
        pixel_data[51][87] = 9;
        pixel_data[51][88] = 10;
        pixel_data[51][89] = 9;
        pixel_data[51][90] = 8;
        pixel_data[51][91] = 6;
        pixel_data[51][92] = 6;
        pixel_data[51][93] = 6;
        pixel_data[51][94] = 4;
        pixel_data[51][95] = 7;
        pixel_data[51][96] = 7;
        pixel_data[51][97] = 12;
        pixel_data[51][98] = 12;
        pixel_data[51][99] = 12; // y=51
        pixel_data[52][0] = 0;
        pixel_data[52][1] = 0;
        pixel_data[52][2] = 0;
        pixel_data[52][3] = 0;
        pixel_data[52][4] = 0;
        pixel_data[52][5] = 6;
        pixel_data[52][6] = 6;
        pixel_data[52][7] = 6;
        pixel_data[52][8] = 6;
        pixel_data[52][9] = 6;
        pixel_data[52][10] = 9;
        pixel_data[52][11] = 10;
        pixel_data[52][12] = 11;
        pixel_data[52][13] = 11;
        pixel_data[52][14] = 11;
        pixel_data[52][15] = 11;
        pixel_data[52][16] = 12;
        pixel_data[52][17] = 12;
        pixel_data[52][18] = 12;
        pixel_data[52][19] = 12;
        pixel_data[52][20] = 12;
        pixel_data[52][21] = 12;
        pixel_data[52][22] = 12;
        pixel_data[52][23] = 12;
        pixel_data[52][24] = 12;
        pixel_data[52][25] = 12;
        pixel_data[52][26] = 13;
        pixel_data[52][27] = 13;
        pixel_data[52][28] = 13;
        pixel_data[52][29] = 13;
        pixel_data[52][30] = 1;
        pixel_data[52][31] = 1;
        pixel_data[52][32] = 13;
        pixel_data[52][33] = 13;
        pixel_data[52][34] = 13;
        pixel_data[52][35] = 13;
        pixel_data[52][36] = 13;
        pixel_data[52][37] = 13;
        pixel_data[52][38] = 1;
        pixel_data[52][39] = 1;
        pixel_data[52][40] = 1;
        pixel_data[52][41] = 13;
        pixel_data[52][42] = 13;
        pixel_data[52][43] = 13;
        pixel_data[52][44] = 13;
        pixel_data[52][45] = 13;
        pixel_data[52][46] = 13;
        pixel_data[52][47] = 13;
        pixel_data[52][48] = 13;
        pixel_data[52][49] = 13;
        pixel_data[52][50] = 13;
        pixel_data[52][51] = 13;
        pixel_data[52][52] = 12;
        pixel_data[52][53] = 12;
        pixel_data[52][54] = 12;
        pixel_data[52][55] = 12;
        pixel_data[52][56] = 12;
        pixel_data[52][57] = 12;
        pixel_data[52][58] = 12;
        pixel_data[52][59] = 12;
        pixel_data[52][60] = 12;
        pixel_data[52][61] = 11;
        pixel_data[52][62] = 11;
        pixel_data[52][63] = 11;
        pixel_data[52][64] = 11;
        pixel_data[52][65] = 11;
        pixel_data[52][66] = 11;
        pixel_data[52][67] = 11;
        pixel_data[52][68] = 11;
        pixel_data[52][69] = 11;
        pixel_data[52][70] = 10;
        pixel_data[52][71] = 10;
        pixel_data[52][72] = 10;
        pixel_data[52][73] = 10;
        pixel_data[52][74] = 10;
        pixel_data[52][75] = 11;
        pixel_data[52][76] = 10;
        pixel_data[52][77] = 10;
        pixel_data[52][78] = 10;
        pixel_data[52][79] = 9;
        pixel_data[52][80] = 8;
        pixel_data[52][81] = 8;
        pixel_data[52][82] = 6;
        pixel_data[52][83] = 6;
        pixel_data[52][84] = 6;
        pixel_data[52][85] = 8;
        pixel_data[52][86] = 8;
        pixel_data[52][87] = 8;
        pixel_data[52][88] = 6;
        pixel_data[52][89] = 6;
        pixel_data[52][90] = 6;
        pixel_data[52][91] = 6;
        pixel_data[52][92] = 8;
        pixel_data[52][93] = 5;
        pixel_data[52][94] = 0;
        pixel_data[52][95] = 0;
        pixel_data[52][96] = 0;
        pixel_data[52][97] = 0;
        pixel_data[52][98] = 0;
        pixel_data[52][99] = 0; // y=52
        pixel_data[53][0] = 0;
        pixel_data[53][1] = 0;
        pixel_data[53][2] = 0;
        pixel_data[53][3] = 0;
        pixel_data[53][4] = 8;
        pixel_data[53][5] = 6;
        pixel_data[53][6] = 6;
        pixel_data[53][7] = 6;
        pixel_data[53][8] = 6;
        pixel_data[53][9] = 6;
        pixel_data[53][10] = 9;
        pixel_data[53][11] = 11;
        pixel_data[53][12] = 11;
        pixel_data[53][13] = 11;
        pixel_data[53][14] = 11;
        pixel_data[53][15] = 11;
        pixel_data[53][16] = 12;
        pixel_data[53][17] = 12;
        pixel_data[53][18] = 12;
        pixel_data[53][19] = 12;
        pixel_data[53][20] = 12;
        pixel_data[53][21] = 12;
        pixel_data[53][22] = 12;
        pixel_data[53][23] = 12;
        pixel_data[53][24] = 12;
        pixel_data[53][25] = 13;
        pixel_data[53][26] = 13;
        pixel_data[53][27] = 13;
        pixel_data[53][28] = 13;
        pixel_data[53][29] = 13;
        pixel_data[53][30] = 13;
        pixel_data[53][31] = 13;
        pixel_data[53][32] = 13;
        pixel_data[53][33] = 13;
        pixel_data[53][34] = 13;
        pixel_data[53][35] = 13;
        pixel_data[53][36] = 13;
        pixel_data[53][37] = 1;
        pixel_data[53][38] = 1;
        pixel_data[53][39] = 1;
        pixel_data[53][40] = 1;
        pixel_data[53][41] = 13;
        pixel_data[53][42] = 13;
        pixel_data[53][43] = 13;
        pixel_data[53][44] = 13;
        pixel_data[53][45] = 13;
        pixel_data[53][46] = 13;
        pixel_data[53][47] = 13;
        pixel_data[53][48] = 13;
        pixel_data[53][49] = 13;
        pixel_data[53][50] = 13;
        pixel_data[53][51] = 13;
        pixel_data[53][52] = 12;
        pixel_data[53][53] = 12;
        pixel_data[53][54] = 12;
        pixel_data[53][55] = 12;
        pixel_data[53][56] = 12;
        pixel_data[53][57] = 12;
        pixel_data[53][58] = 12;
        pixel_data[53][59] = 12;
        pixel_data[53][60] = 12;
        pixel_data[53][61] = 11;
        pixel_data[53][62] = 11;
        pixel_data[53][63] = 11;
        pixel_data[53][64] = 11;
        pixel_data[53][65] = 11;
        pixel_data[53][66] = 11;
        pixel_data[53][67] = 11;
        pixel_data[53][68] = 11;
        pixel_data[53][69] = 10;
        pixel_data[53][70] = 10;
        pixel_data[53][71] = 10;
        pixel_data[53][72] = 10;
        pixel_data[53][73] = 10;
        pixel_data[53][74] = 11;
        pixel_data[53][75] = 10;
        pixel_data[53][76] = 10;
        pixel_data[53][77] = 9;
        pixel_data[53][78] = 8;
        pixel_data[53][79] = 6;
        pixel_data[53][80] = 6;
        pixel_data[53][81] = 6;
        pixel_data[53][82] = 6;
        pixel_data[53][83] = 6;
        pixel_data[53][84] = 6;
        pixel_data[53][85] = 6;
        pixel_data[53][86] = 6;
        pixel_data[53][87] = 6;
        pixel_data[53][88] = 6;
        pixel_data[53][89] = 6;
        pixel_data[53][90] = 6;
        pixel_data[53][91] = 5;
        pixel_data[53][92] = 7;
        pixel_data[53][93] = 0;
        pixel_data[53][94] = 0;
        pixel_data[53][95] = 0;
        pixel_data[53][96] = 0;
        pixel_data[53][97] = 0;
        pixel_data[53][98] = 0;
        pixel_data[53][99] = 0; // y=53
        pixel_data[54][0] = 0;
        pixel_data[54][1] = 0;
        pixel_data[54][2] = 0;
        pixel_data[54][3] = 5;
        pixel_data[54][4] = 6;
        pixel_data[54][5] = 6;
        pixel_data[54][6] = 6;
        pixel_data[54][7] = 6;
        pixel_data[54][8] = 6;
        pixel_data[54][9] = 8;
        pixel_data[54][10] = 9;
        pixel_data[54][11] = 10;
        pixel_data[54][12] = 11;
        pixel_data[54][13] = 11;
        pixel_data[54][14] = 11;
        pixel_data[54][15] = 11;
        pixel_data[54][16] = 12;
        pixel_data[54][17] = 12;
        pixel_data[54][18] = 12;
        pixel_data[54][19] = 12;
        pixel_data[54][20] = 12;
        pixel_data[54][21] = 12;
        pixel_data[54][22] = 12;
        pixel_data[54][23] = 12;
        pixel_data[54][24] = 13;
        pixel_data[54][25] = 13;
        pixel_data[54][26] = 13;
        pixel_data[54][27] = 13;
        pixel_data[54][28] = 13;
        pixel_data[54][29] = 13;
        pixel_data[54][30] = 13;
        pixel_data[54][31] = 13;
        pixel_data[54][32] = 13;
        pixel_data[54][33] = 13;
        pixel_data[54][34] = 13;
        pixel_data[54][35] = 13;
        pixel_data[54][36] = 13;
        pixel_data[54][37] = 1;
        pixel_data[54][38] = 1;
        pixel_data[54][39] = 1;
        pixel_data[54][40] = 13;
        pixel_data[54][41] = 13;
        pixel_data[54][42] = 13;
        pixel_data[54][43] = 13;
        pixel_data[54][44] = 13;
        pixel_data[54][45] = 13;
        pixel_data[54][46] = 13;
        pixel_data[54][47] = 13;
        pixel_data[54][48] = 13;
        pixel_data[54][49] = 13;
        pixel_data[54][50] = 13;
        pixel_data[54][51] = 12;
        pixel_data[54][52] = 12;
        pixel_data[54][53] = 12;
        pixel_data[54][54] = 12;
        pixel_data[54][55] = 12;
        pixel_data[54][56] = 12;
        pixel_data[54][57] = 12;
        pixel_data[54][58] = 12;
        pixel_data[54][59] = 12;
        pixel_data[54][60] = 12;
        pixel_data[54][61] = 11;
        pixel_data[54][62] = 11;
        pixel_data[54][63] = 11;
        pixel_data[54][64] = 11;
        pixel_data[54][65] = 11;
        pixel_data[54][66] = 11;
        pixel_data[54][67] = 11;
        pixel_data[54][68] = 11;
        pixel_data[54][69] = 11;
        pixel_data[54][70] = 11;
        pixel_data[54][71] = 10;
        pixel_data[54][72] = 10;
        pixel_data[54][73] = 10;
        pixel_data[54][74] = 10;
        pixel_data[54][75] = 9;
        pixel_data[54][76] = 8;
        pixel_data[54][77] = 6;
        pixel_data[54][78] = 4;
        pixel_data[54][79] = 4;
        pixel_data[54][80] = 6;
        pixel_data[54][81] = 6;
        pixel_data[54][82] = 6;
        pixel_data[54][83] = 6;
        pixel_data[54][84] = 6;
        pixel_data[54][85] = 6;
        pixel_data[54][86] = 6;
        pixel_data[54][87] = 6;
        pixel_data[54][88] = 6;
        pixel_data[54][89] = 6;
        pixel_data[54][90] = 6;
        pixel_data[54][91] = 6;
        pixel_data[54][92] = 0;
        pixel_data[54][93] = 0;
        pixel_data[54][94] = 0;
        pixel_data[54][95] = 0;
        pixel_data[54][96] = 0;
        pixel_data[54][97] = 0;
        pixel_data[54][98] = 0;
        pixel_data[54][99] = 0; // y=54
        pixel_data[55][0] = 0;
        pixel_data[55][1] = 0;
        pixel_data[55][2] = 1;
        pixel_data[55][3] = 5;
        pixel_data[55][4] = 6;
        pixel_data[55][5] = 6;
        pixel_data[55][6] = 6;
        pixel_data[55][7] = 6;
        pixel_data[55][8] = 6;
        pixel_data[55][9] = 6;
        pixel_data[55][10] = 9;
        pixel_data[55][11] = 10;
        pixel_data[55][12] = 11;
        pixel_data[55][13] = 11;
        pixel_data[55][14] = 11;
        pixel_data[55][15] = 11;
        pixel_data[55][16] = 12;
        pixel_data[55][17] = 12;
        pixel_data[55][18] = 12;
        pixel_data[55][19] = 12;
        pixel_data[55][20] = 12;
        pixel_data[55][21] = 12;
        pixel_data[55][22] = 12;
        pixel_data[55][23] = 12;
        pixel_data[55][24] = 13;
        pixel_data[55][25] = 13;
        pixel_data[55][26] = 13;
        pixel_data[55][27] = 13;
        pixel_data[55][28] = 13;
        pixel_data[55][29] = 13;
        pixel_data[55][30] = 13;
        pixel_data[55][31] = 13;
        pixel_data[55][32] = 13;
        pixel_data[55][33] = 13;
        pixel_data[55][34] = 13;
        pixel_data[55][35] = 13;
        pixel_data[55][36] = 1;
        pixel_data[55][37] = 1;
        pixel_data[55][38] = 1;
        pixel_data[55][39] = 1;
        pixel_data[55][40] = 13;
        pixel_data[55][41] = 13;
        pixel_data[55][42] = 13;
        pixel_data[55][43] = 13;
        pixel_data[55][44] = 13;
        pixel_data[55][45] = 13;
        pixel_data[55][46] = 13;
        pixel_data[55][47] = 13;
        pixel_data[55][48] = 13;
        pixel_data[55][49] = 13;
        pixel_data[55][50] = 12;
        pixel_data[55][51] = 12;
        pixel_data[55][52] = 12;
        pixel_data[55][53] = 12;
        pixel_data[55][54] = 12;
        pixel_data[55][55] = 12;
        pixel_data[55][56] = 12;
        pixel_data[55][57] = 12;
        pixel_data[55][58] = 12;
        pixel_data[55][59] = 12;
        pixel_data[55][60] = 11;
        pixel_data[55][61] = 11;
        pixel_data[55][62] = 11;
        pixel_data[55][63] = 11;
        pixel_data[55][64] = 11;
        pixel_data[55][65] = 11;
        pixel_data[55][66] = 11;
        pixel_data[55][67] = 11;
        pixel_data[55][68] = 11;
        pixel_data[55][69] = 11;
        pixel_data[55][70] = 10;
        pixel_data[55][71] = 10;
        pixel_data[55][72] = 9;
        pixel_data[55][73] = 8;
        pixel_data[55][74] = 6;
        pixel_data[55][75] = 4;
        pixel_data[55][76] = 4;
        pixel_data[55][77] = 4;
        pixel_data[55][78] = 4;
        pixel_data[55][79] = 6;
        pixel_data[55][80] = 6;
        pixel_data[55][81] = 6;
        pixel_data[55][82] = 6;
        pixel_data[55][83] = 6;
        pixel_data[55][84] = 6;
        pixel_data[55][85] = 6;
        pixel_data[55][86] = 6;
        pixel_data[55][87] = 6;
        pixel_data[55][88] = 6;
        pixel_data[55][89] = 6;
        pixel_data[55][90] = 7;
        pixel_data[55][91] = 0;
        pixel_data[55][92] = 0;
        pixel_data[55][93] = 0;
        pixel_data[55][94] = 0;
        pixel_data[55][95] = 0;
        pixel_data[55][96] = 0;
        pixel_data[55][97] = 0;
        pixel_data[55][98] = 0;
        pixel_data[55][99] = 0; // y=55
        pixel_data[56][0] = 0;
        pixel_data[56][1] = 0;
        pixel_data[56][2] = 1;
        pixel_data[56][3] = 8;
        pixel_data[56][4] = 6;
        pixel_data[56][5] = 6;
        pixel_data[56][6] = 6;
        pixel_data[56][7] = 6;
        pixel_data[56][8] = 6;
        pixel_data[56][9] = 6;
        pixel_data[56][10] = 8;
        pixel_data[56][11] = 10;
        pixel_data[56][12] = 11;
        pixel_data[56][13] = 11;
        pixel_data[56][14] = 11;
        pixel_data[56][15] = 11;
        pixel_data[56][16] = 12;
        pixel_data[56][17] = 12;
        pixel_data[56][18] = 12;
        pixel_data[56][19] = 12;
        pixel_data[56][20] = 12;
        pixel_data[56][21] = 12;
        pixel_data[56][22] = 12;
        pixel_data[56][23] = 12;
        pixel_data[56][24] = 13;
        pixel_data[56][25] = 13;
        pixel_data[56][26] = 13;
        pixel_data[56][27] = 13;
        pixel_data[56][28] = 13;
        pixel_data[56][29] = 13;
        pixel_data[56][30] = 13;
        pixel_data[56][31] = 13;
        pixel_data[56][32] = 13;
        pixel_data[56][33] = 13;
        pixel_data[56][34] = 13;
        pixel_data[56][35] = 1;
        pixel_data[56][36] = 1;
        pixel_data[56][37] = 1;
        pixel_data[56][38] = 1;
        pixel_data[56][39] = 1;
        pixel_data[56][40] = 13;
        pixel_data[56][41] = 13;
        pixel_data[56][42] = 13;
        pixel_data[56][43] = 13;
        pixel_data[56][44] = 13;
        pixel_data[56][45] = 13;
        pixel_data[56][46] = 13;
        pixel_data[56][47] = 13;
        pixel_data[56][48] = 13;
        pixel_data[56][49] = 13;
        pixel_data[56][50] = 12;
        pixel_data[56][51] = 12;
        pixel_data[56][52] = 12;
        pixel_data[56][53] = 12;
        pixel_data[56][54] = 12;
        pixel_data[56][55] = 12;
        pixel_data[56][56] = 12;
        pixel_data[56][57] = 12;
        pixel_data[56][58] = 12;
        pixel_data[56][59] = 11;
        pixel_data[56][60] = 11;
        pixel_data[56][61] = 11;
        pixel_data[56][62] = 11;
        pixel_data[56][63] = 11;
        pixel_data[56][64] = 11;
        pixel_data[56][65] = 11;
        pixel_data[56][66] = 11;
        pixel_data[56][67] = 10;
        pixel_data[56][68] = 10;
        pixel_data[56][69] = 9;
        pixel_data[56][70] = 8;
        pixel_data[56][71] = 6;
        pixel_data[56][72] = 4;
        pixel_data[56][73] = 4;
        pixel_data[56][74] = 4;
        pixel_data[56][75] = 4;
        pixel_data[56][76] = 6;
        pixel_data[56][77] = 6;
        pixel_data[56][78] = 6;
        pixel_data[56][79] = 6;
        pixel_data[56][80] = 6;
        pixel_data[56][81] = 6;
        pixel_data[56][82] = 6;
        pixel_data[56][83] = 6;
        pixel_data[56][84] = 6;
        pixel_data[56][85] = 6;
        pixel_data[56][86] = 6;
        pixel_data[56][87] = 6;
        pixel_data[56][88] = 8;
        pixel_data[56][89] = 14;
        pixel_data[56][90] = 0;
        pixel_data[56][91] = 0;
        pixel_data[56][92] = 0;
        pixel_data[56][93] = 0;
        pixel_data[56][94] = 0;
        pixel_data[56][95] = 0;
        pixel_data[56][96] = 0;
        pixel_data[56][97] = 0;
        pixel_data[56][98] = 0;
        pixel_data[56][99] = 0; // y=56
        pixel_data[57][0] = 0;
        pixel_data[57][1] = 0;
        pixel_data[57][2] = 1;
        pixel_data[57][3] = 8;
        pixel_data[57][4] = 6;
        pixel_data[57][5] = 6;
        pixel_data[57][6] = 6;
        pixel_data[57][7] = 6;
        pixel_data[57][8] = 6;
        pixel_data[57][9] = 6;
        pixel_data[57][10] = 8;
        pixel_data[57][11] = 9;
        pixel_data[57][12] = 10;
        pixel_data[57][13] = 10;
        pixel_data[57][14] = 11;
        pixel_data[57][15] = 11;
        pixel_data[57][16] = 11;
        pixel_data[57][17] = 12;
        pixel_data[57][18] = 12;
        pixel_data[57][19] = 12;
        pixel_data[57][20] = 12;
        pixel_data[57][21] = 12;
        pixel_data[57][22] = 12;
        pixel_data[57][23] = 12;
        pixel_data[57][24] = 12;
        pixel_data[57][25] = 13;
        pixel_data[57][26] = 13;
        pixel_data[57][27] = 13;
        pixel_data[57][28] = 13;
        pixel_data[57][29] = 13;
        pixel_data[57][30] = 13;
        pixel_data[57][31] = 13;
        pixel_data[57][32] = 13;
        pixel_data[57][33] = 13;
        pixel_data[57][34] = 13;
        pixel_data[57][35] = 1;
        pixel_data[57][36] = 1;
        pixel_data[57][37] = 1;
        pixel_data[57][38] = 1;
        pixel_data[57][39] = 1;
        pixel_data[57][40] = 13;
        pixel_data[57][41] = 13;
        pixel_data[57][42] = 13;
        pixel_data[57][43] = 13;
        pixel_data[57][44] = 13;
        pixel_data[57][45] = 13;
        pixel_data[57][46] = 13;
        pixel_data[57][47] = 13;
        pixel_data[57][48] = 13;
        pixel_data[57][49] = 12;
        pixel_data[57][50] = 12;
        pixel_data[57][51] = 12;
        pixel_data[57][52] = 12;
        pixel_data[57][53] = 12;
        pixel_data[57][54] = 12;
        pixel_data[57][55] = 12;
        pixel_data[57][56] = 12;
        pixel_data[57][57] = 12;
        pixel_data[57][58] = 12;
        pixel_data[57][59] = 12;
        pixel_data[57][60] = 12;
        pixel_data[57][61] = 11;
        pixel_data[57][62] = 11;
        pixel_data[57][63] = 11;
        pixel_data[57][64] = 10;
        pixel_data[57][65] = 10;
        pixel_data[57][66] = 9;
        pixel_data[57][67] = 8;
        pixel_data[57][68] = 6;
        pixel_data[57][69] = 4;
        pixel_data[57][70] = 4;
        pixel_data[57][71] = 4;
        pixel_data[57][72] = 4;
        pixel_data[57][73] = 4;
        pixel_data[57][74] = 6;
        pixel_data[57][75] = 6;
        pixel_data[57][76] = 6;
        pixel_data[57][77] = 6;
        pixel_data[57][78] = 6;
        pixel_data[57][79] = 6;
        pixel_data[57][80] = 6;
        pixel_data[57][81] = 6;
        pixel_data[57][82] = 4;
        pixel_data[57][83] = 6;
        pixel_data[57][84] = 7;
        pixel_data[57][85] = 2;
        pixel_data[57][86] = 7;
        pixel_data[57][87] = 1;
        pixel_data[57][88] = 0;
        pixel_data[57][89] = 0;
        pixel_data[57][90] = 0;
        pixel_data[57][91] = 0;
        pixel_data[57][92] = 0;
        pixel_data[57][93] = 0;
        pixel_data[57][94] = 0;
        pixel_data[57][95] = 0;
        pixel_data[57][96] = 0;
        pixel_data[57][97] = 0;
        pixel_data[57][98] = 0;
        pixel_data[57][99] = 0; // y=57
        pixel_data[58][0] = 0;
        pixel_data[58][1] = 0;
        pixel_data[58][2] = 0;
        pixel_data[58][3] = 7;
        pixel_data[58][4] = 6;
        pixel_data[58][5] = 6;
        pixel_data[58][6] = 6;
        pixel_data[58][7] = 6;
        pixel_data[58][8] = 6;
        pixel_data[58][9] = 6;
        pixel_data[58][10] = 6;
        pixel_data[58][11] = 6;
        pixel_data[58][12] = 9;
        pixel_data[58][13] = 9;
        pixel_data[58][14] = 10;
        pixel_data[58][15] = 10;
        pixel_data[58][16] = 11;
        pixel_data[58][17] = 11;
        pixel_data[58][18] = 12;
        pixel_data[58][19] = 12;
        pixel_data[58][20] = 12;
        pixel_data[58][21] = 12;
        pixel_data[58][22] = 12;
        pixel_data[58][23] = 12;
        pixel_data[58][24] = 12;
        pixel_data[58][25] = 12;
        pixel_data[58][26] = 12;
        pixel_data[58][27] = 12;
        pixel_data[58][28] = 12;
        pixel_data[58][29] = 13;
        pixel_data[58][30] = 13;
        pixel_data[58][31] = 13;
        pixel_data[58][32] = 13;
        pixel_data[58][33] = 13;
        pixel_data[58][34] = 1;
        pixel_data[58][35] = 1;
        pixel_data[58][36] = 1;
        pixel_data[58][37] = 1;
        pixel_data[58][38] = 1;
        pixel_data[58][39] = 1;
        pixel_data[58][40] = 13;
        pixel_data[58][41] = 13;
        pixel_data[58][42] = 13;
        pixel_data[58][43] = 13;
        pixel_data[58][44] = 13;
        pixel_data[58][45] = 13;
        pixel_data[58][46] = 13;
        pixel_data[58][47] = 13;
        pixel_data[58][48] = 12;
        pixel_data[58][49] = 12;
        pixel_data[58][50] = 12;
        pixel_data[58][51] = 12;
        pixel_data[58][52] = 12;
        pixel_data[58][53] = 12;
        pixel_data[58][54] = 12;
        pixel_data[58][55] = 12;
        pixel_data[58][56] = 12;
        pixel_data[58][57] = 12;
        pixel_data[58][58] = 12;
        pixel_data[58][59] = 11;
        pixel_data[58][60] = 11;
        pixel_data[58][61] = 10;
        pixel_data[58][62] = 10;
        pixel_data[58][63] = 9;
        pixel_data[58][64] = 6;
        pixel_data[58][65] = 6;
        pixel_data[58][66] = 4;
        pixel_data[58][67] = 4;
        pixel_data[58][68] = 4;
        pixel_data[58][69] = 4;
        pixel_data[58][70] = 6;
        pixel_data[58][71] = 6;
        pixel_data[58][72] = 6;
        pixel_data[58][73] = 6;
        pixel_data[58][74] = 6;
        pixel_data[58][75] = 6;
        pixel_data[58][76] = 6;
        pixel_data[58][77] = 6;
        pixel_data[58][78] = 6;
        pixel_data[58][79] = 5;
        pixel_data[58][80] = 7;
        pixel_data[58][81] = 2;
        pixel_data[58][82] = 1;
        pixel_data[58][83] = 0;
        pixel_data[58][84] = 0;
        pixel_data[58][85] = 0;
        pixel_data[58][86] = 0;
        pixel_data[58][87] = 0;
        pixel_data[58][88] = 0;
        pixel_data[58][89] = 0;
        pixel_data[58][90] = 0;
        pixel_data[58][91] = 0;
        pixel_data[58][92] = 0;
        pixel_data[58][93] = 0;
        pixel_data[58][94] = 0;
        pixel_data[58][95] = 0;
        pixel_data[58][96] = 0;
        pixel_data[58][97] = 0;
        pixel_data[58][98] = 0;
        pixel_data[58][99] = 0; // y=58
        pixel_data[59][0] = 0;
        pixel_data[59][1] = 0;
        pixel_data[59][2] = 0;
        pixel_data[59][3] = 1;
        pixel_data[59][4] = 6;
        pixel_data[59][5] = 6;
        pixel_data[59][6] = 6;
        pixel_data[59][7] = 6;
        pixel_data[59][8] = 6;
        pixel_data[59][9] = 6;
        pixel_data[59][10] = 6;
        pixel_data[59][11] = 6;
        pixel_data[59][12] = 6;
        pixel_data[59][13] = 8;
        pixel_data[59][14] = 9;
        pixel_data[59][15] = 10;
        pixel_data[59][16] = 11;
        pixel_data[59][17] = 11;
        pixel_data[59][18] = 12;
        pixel_data[59][19] = 12;
        pixel_data[59][20] = 12;
        pixel_data[59][21] = 12;
        pixel_data[59][22] = 12;
        pixel_data[59][23] = 12;
        pixel_data[59][24] = 12;
        pixel_data[59][25] = 12;
        pixel_data[59][26] = 12;
        pixel_data[59][27] = 12;
        pixel_data[59][28] = 12;
        pixel_data[59][29] = 12;
        pixel_data[59][30] = 13;
        pixel_data[59][31] = 13;
        pixel_data[59][32] = 13;
        pixel_data[59][33] = 1;
        pixel_data[59][34] = 1;
        pixel_data[59][35] = 1;
        pixel_data[59][36] = 1;
        pixel_data[59][37] = 1;
        pixel_data[59][38] = 1;
        pixel_data[59][39] = 1;
        pixel_data[59][40] = 13;
        pixel_data[59][41] = 13;
        pixel_data[59][42] = 13;
        pixel_data[59][43] = 13;
        pixel_data[59][44] = 13;
        pixel_data[59][45] = 13;
        pixel_data[59][46] = 13;
        pixel_data[59][47] = 13;
        pixel_data[59][48] = 13;
        pixel_data[59][49] = 13;
        pixel_data[59][50] = 13;
        pixel_data[59][51] = 12;
        pixel_data[59][52] = 12;
        pixel_data[59][53] = 12;
        pixel_data[59][54] = 12;
        pixel_data[59][55] = 12;
        pixel_data[59][56] = 11;
        pixel_data[59][57] = 11;
        pixel_data[59][58] = 10;
        pixel_data[59][59] = 9;
        pixel_data[59][60] = 9;
        pixel_data[59][61] = 8;
        pixel_data[59][62] = 6;
        pixel_data[59][63] = 6;
        pixel_data[59][64] = 4;
        pixel_data[59][65] = 4;
        pixel_data[59][66] = 4;
        pixel_data[59][67] = 6;
        pixel_data[59][68] = 6;
        pixel_data[59][69] = 6;
        pixel_data[59][70] = 6;
        pixel_data[59][71] = 6;
        pixel_data[59][72] = 6;
        pixel_data[59][73] = 6;
        pixel_data[59][74] = 6;
        pixel_data[59][75] = 6;
        pixel_data[59][76] = 6;
        pixel_data[59][77] = 6;
        pixel_data[59][78] = 2;
        pixel_data[59][79] = 0;
        pixel_data[59][80] = 0;
        pixel_data[59][81] = 0;
        pixel_data[59][82] = 0;
        pixel_data[59][83] = 0;
        pixel_data[59][84] = 0;
        pixel_data[59][85] = 0;
        pixel_data[59][86] = 0;
        pixel_data[59][87] = 0;
        pixel_data[59][88] = 0;
        pixel_data[59][89] = 0;
        pixel_data[59][90] = 0;
        pixel_data[59][91] = 0;
        pixel_data[59][92] = 0;
        pixel_data[59][93] = 0;
        pixel_data[59][94] = 0;
        pixel_data[59][95] = 0;
        pixel_data[59][96] = 0;
        pixel_data[59][97] = 0;
        pixel_data[59][98] = 0;
        pixel_data[59][99] = 0; // y=59
        pixel_data[60][0] = 0;
        pixel_data[60][1] = 0;
        pixel_data[60][2] = 0;
        pixel_data[60][3] = 0;
        pixel_data[60][4] = 7;
        pixel_data[60][5] = 6;
        pixel_data[60][6] = 6;
        pixel_data[60][7] = 6;
        pixel_data[60][8] = 6;
        pixel_data[60][9] = 6;
        pixel_data[60][10] = 6;
        pixel_data[60][11] = 5;
        pixel_data[60][12] = 8;
        pixel_data[60][13] = 6;
        pixel_data[60][14] = 9;
        pixel_data[60][15] = 10;
        pixel_data[60][16] = 11;
        pixel_data[60][17] = 12;
        pixel_data[60][18] = 12;
        pixel_data[60][19] = 12;
        pixel_data[60][20] = 12;
        pixel_data[60][21] = 12;
        pixel_data[60][22] = 12;
        pixel_data[60][23] = 12;
        pixel_data[60][24] = 12;
        pixel_data[60][25] = 12;
        pixel_data[60][26] = 12;
        pixel_data[60][27] = 12;
        pixel_data[60][28] = 12;
        pixel_data[60][29] = 12;
        pixel_data[60][30] = 12;
        pixel_data[60][31] = 13;
        pixel_data[60][32] = 13;
        pixel_data[60][33] = 1;
        pixel_data[60][34] = 1;
        pixel_data[60][35] = 1;
        pixel_data[60][36] = 1;
        pixel_data[60][37] = 1;
        pixel_data[60][38] = 1;
        pixel_data[60][39] = 1;
        pixel_data[60][40] = 1;
        pixel_data[60][41] = 13;
        pixel_data[60][42] = 13;
        pixel_data[60][43] = 13;
        pixel_data[60][44] = 13;
        pixel_data[60][45] = 13;
        pixel_data[60][46] = 13;
        pixel_data[60][47] = 13;
        pixel_data[60][48] = 13;
        pixel_data[60][49] = 13;
        pixel_data[60][50] = 13;
        pixel_data[60][51] = 12;
        pixel_data[60][52] = 11;
        pixel_data[60][53] = 11;
        pixel_data[60][54] = 10;
        pixel_data[60][55] = 10;
        pixel_data[60][56] = 9;
        pixel_data[60][57] = 9;
        pixel_data[60][58] = 8;
        pixel_data[60][59] = 8;
        pixel_data[60][60] = 6;
        pixel_data[60][61] = 6;
        pixel_data[60][62] = 6;
        pixel_data[60][63] = 6;
        pixel_data[60][64] = 6;
        pixel_data[60][65] = 6;
        pixel_data[60][66] = 6;
        pixel_data[60][67] = 6;
        pixel_data[60][68] = 6;
        pixel_data[60][69] = 6;
        pixel_data[60][70] = 6;
        pixel_data[60][71] = 6;
        pixel_data[60][72] = 6;
        pixel_data[60][73] = 6;
        pixel_data[60][74] = 6;
        pixel_data[60][75] = 10;
        pixel_data[60][76] = 1;
        pixel_data[60][77] = 0;
        pixel_data[60][78] = 0;
        pixel_data[60][79] = 0;
        pixel_data[60][80] = 0;
        pixel_data[60][81] = 0;
        pixel_data[60][82] = 0;
        pixel_data[60][83] = 0;
        pixel_data[60][84] = 0;
        pixel_data[60][85] = 0;
        pixel_data[60][86] = 0;
        pixel_data[60][87] = 0;
        pixel_data[60][88] = 0;
        pixel_data[60][89] = 0;
        pixel_data[60][90] = 0;
        pixel_data[60][91] = 0;
        pixel_data[60][92] = 0;
        pixel_data[60][93] = 0;
        pixel_data[60][94] = 0;
        pixel_data[60][95] = 0;
        pixel_data[60][96] = 0;
        pixel_data[60][97] = 0;
        pixel_data[60][98] = 0;
        pixel_data[60][99] = 0; // y=60
        pixel_data[61][0] = 0;
        pixel_data[61][1] = 0;
        pixel_data[61][2] = 0;
        pixel_data[61][3] = 0;
        pixel_data[61][4] = 0;
        pixel_data[61][5] = 7;
        pixel_data[61][6] = 15;
        pixel_data[61][7] = 2;
        pixel_data[61][8] = 7;
        pixel_data[61][9] = 2;
        pixel_data[61][10] = 15;
        pixel_data[61][11] = 7;
        pixel_data[61][12] = 6;
        pixel_data[61][13] = 8;
        pixel_data[61][14] = 9;
        pixel_data[61][15] = 10;
        pixel_data[61][16] = 11;
        pixel_data[61][17] = 12;
        pixel_data[61][18] = 12;
        pixel_data[61][19] = 12;
        pixel_data[61][20] = 12;
        pixel_data[61][21] = 12;
        pixel_data[61][22] = 12;
        pixel_data[61][23] = 12;
        pixel_data[61][24] = 12;
        pixel_data[61][25] = 12;
        pixel_data[61][26] = 12;
        pixel_data[61][27] = 12;
        pixel_data[61][28] = 12;
        pixel_data[61][29] = 12;
        pixel_data[61][30] = 12;
        pixel_data[61][31] = 12;
        pixel_data[61][32] = 13;
        pixel_data[61][33] = 13;
        pixel_data[61][34] = 1;
        pixel_data[61][35] = 1;
        pixel_data[61][36] = 1;
        pixel_data[61][37] = 1;
        pixel_data[61][38] = 1;
        pixel_data[61][39] = 1;
        pixel_data[61][40] = 1;
        pixel_data[61][41] = 1;
        pixel_data[61][42] = 13;
        pixel_data[61][43] = 13;
        pixel_data[61][44] = 12;
        pixel_data[61][45] = 12;
        pixel_data[61][46] = 12;
        pixel_data[61][47] = 11;
        pixel_data[61][48] = 11;
        pixel_data[61][49] = 10;
        pixel_data[61][50] = 10;
        pixel_data[61][51] = 9;
        pixel_data[61][52] = 9;
        pixel_data[61][53] = 9;
        pixel_data[61][54] = 9;
        pixel_data[61][55] = 9;
        pixel_data[61][56] = 8;
        pixel_data[61][57] = 6;
        pixel_data[61][58] = 6;
        pixel_data[61][59] = 6;
        pixel_data[61][60] = 6;
        pixel_data[61][61] = 6;
        pixel_data[61][62] = 6;
        pixel_data[61][63] = 6;
        pixel_data[61][64] = 6;
        pixel_data[61][65] = 6;
        pixel_data[61][66] = 6;
        pixel_data[61][67] = 6;
        pixel_data[61][68] = 6;
        pixel_data[61][69] = 6;
        pixel_data[61][70] = 6;
        pixel_data[61][71] = 6;
        pixel_data[61][72] = 6;
        pixel_data[61][73] = 7;
        pixel_data[61][74] = 15;
        pixel_data[61][75] = 0;
        pixel_data[61][76] = 0;
        pixel_data[61][77] = 0;
        pixel_data[61][78] = 0;
        pixel_data[61][79] = 0;
        pixel_data[61][80] = 0;
        pixel_data[61][81] = 0;
        pixel_data[61][82] = 0;
        pixel_data[61][83] = 0;
        pixel_data[61][84] = 0;
        pixel_data[61][85] = 0;
        pixel_data[61][86] = 0;
        pixel_data[61][87] = 0;
        pixel_data[61][88] = 0;
        pixel_data[61][89] = 0;
        pixel_data[61][90] = 0;
        pixel_data[61][91] = 0;
        pixel_data[61][92] = 0;
        pixel_data[61][93] = 0;
        pixel_data[61][94] = 0;
        pixel_data[61][95] = 0;
        pixel_data[61][96] = 0;
        pixel_data[61][97] = 0;
        pixel_data[61][98] = 0;
        pixel_data[61][99] = 0; // y=61
        pixel_data[62][0] = 0;
        pixel_data[62][1] = 0;
        pixel_data[62][2] = 0;
        pixel_data[62][3] = 0;
        pixel_data[62][4] = 0;
        pixel_data[62][5] = 0;
        pixel_data[62][6] = 0;
        pixel_data[62][7] = 0;
        pixel_data[62][8] = 0;
        pixel_data[62][9] = 0;
        pixel_data[62][10] = 0;
        pixel_data[62][11] = 5;
        pixel_data[62][12] = 6;
        pixel_data[62][13] = 8;
        pixel_data[62][14] = 10;
        pixel_data[62][15] = 11;
        pixel_data[62][16] = 11;
        pixel_data[62][17] = 11;
        pixel_data[62][18] = 11;
        pixel_data[62][19] = 12;
        pixel_data[62][20] = 12;
        pixel_data[62][21] = 12;
        pixel_data[62][22] = 12;
        pixel_data[62][23] = 12;
        pixel_data[62][24] = 12;
        pixel_data[62][25] = 12;
        pixel_data[62][26] = 12;
        pixel_data[62][27] = 12;
        pixel_data[62][28] = 12;
        pixel_data[62][29] = 11;
        pixel_data[62][30] = 11;
        pixel_data[62][31] = 11;
        pixel_data[62][32] = 11;
        pixel_data[62][33] = 11;
        pixel_data[62][34] = 12;
        pixel_data[62][35] = 12;
        pixel_data[62][36] = 12;
        pixel_data[62][37] = 12;
        pixel_data[62][38] = 12;
        pixel_data[62][39] = 11;
        pixel_data[62][40] = 11;
        pixel_data[62][41] = 11;
        pixel_data[62][42] = 10;
        pixel_data[62][43] = 10;
        pixel_data[62][44] = 10;
        pixel_data[62][45] = 9;
        pixel_data[62][46] = 9;
        pixel_data[62][47] = 8;
        pixel_data[62][48] = 8;
        pixel_data[62][49] = 8;
        pixel_data[62][50] = 8;
        pixel_data[62][51] = 8;
        pixel_data[62][52] = 8;
        pixel_data[62][53] = 8;
        pixel_data[62][54] = 8;
        pixel_data[62][55] = 6;
        pixel_data[62][56] = 6;
        pixel_data[62][57] = 6;
        pixel_data[62][58] = 6;
        pixel_data[62][59] = 6;
        pixel_data[62][60] = 6;
        pixel_data[62][61] = 6;
        pixel_data[62][62] = 6;
        pixel_data[62][63] = 6;
        pixel_data[62][64] = 6;
        pixel_data[62][65] = 6;
        pixel_data[62][66] = 6;
        pixel_data[62][67] = 6;
        pixel_data[62][68] = 6;
        pixel_data[62][69] = 6;
        pixel_data[62][70] = 6;
        pixel_data[62][71] = 8;
        pixel_data[62][72] = 7;
        pixel_data[62][73] = 0;
        pixel_data[62][74] = 0;
        pixel_data[62][75] = 0;
        pixel_data[62][76] = 0;
        pixel_data[62][77] = 0;
        pixel_data[62][78] = 0;
        pixel_data[62][79] = 0;
        pixel_data[62][80] = 0;
        pixel_data[62][81] = 0;
        pixel_data[62][82] = 0;
        pixel_data[62][83] = 0;
        pixel_data[62][84] = 0;
        pixel_data[62][85] = 0;
        pixel_data[62][86] = 0;
        pixel_data[62][87] = 0;
        pixel_data[62][88] = 0;
        pixel_data[62][89] = 0;
        pixel_data[62][90] = 0;
        pixel_data[62][91] = 0;
        pixel_data[62][92] = 0;
        pixel_data[62][93] = 0;
        pixel_data[62][94] = 0;
        pixel_data[62][95] = 0;
        pixel_data[62][96] = 0;
        pixel_data[62][97] = 0;
        pixel_data[62][98] = 0;
        pixel_data[62][99] = 0; // y=62
        pixel_data[63][0] = 0;
        pixel_data[63][1] = 0;
        pixel_data[63][2] = 0;
        pixel_data[63][3] = 0;
        pixel_data[63][4] = 0;
        pixel_data[63][5] = 0;
        pixel_data[63][6] = 0;
        pixel_data[63][7] = 0;
        pixel_data[63][8] = 0;
        pixel_data[63][9] = 0;
        pixel_data[63][10] = 0;
        pixel_data[63][11] = 9;
        pixel_data[63][12] = 8;
        pixel_data[63][13] = 9;
        pixel_data[63][14] = 10;
        pixel_data[63][15] = 11;
        pixel_data[63][16] = 11;
        pixel_data[63][17] = 11;
        pixel_data[63][18] = 11;
        pixel_data[63][19] = 11;
        pixel_data[63][20] = 12;
        pixel_data[63][21] = 12;
        pixel_data[63][22] = 12;
        pixel_data[63][23] = 12;
        pixel_data[63][24] = 12;
        pixel_data[63][25] = 12;
        pixel_data[63][26] = 12;
        pixel_data[63][27] = 12;
        pixel_data[63][28] = 12;
        pixel_data[63][29] = 11;
        pixel_data[63][30] = 11;
        pixel_data[63][31] = 10;
        pixel_data[63][32] = 10;
        pixel_data[63][33] = 10;
        pixel_data[63][34] = 10;
        pixel_data[63][35] = 9;
        pixel_data[63][36] = 9;
        pixel_data[63][37] = 9;
        pixel_data[63][38] = 8;
        pixel_data[63][39] = 8;
        pixel_data[63][40] = 8;
        pixel_data[63][41] = 8;
        pixel_data[63][42] = 8;
        pixel_data[63][43] = 6;
        pixel_data[63][44] = 6;
        pixel_data[63][45] = 6;
        pixel_data[63][46] = 6;
        pixel_data[63][47] = 6;
        pixel_data[63][48] = 6;
        pixel_data[63][49] = 6;
        pixel_data[63][50] = 6;
        pixel_data[63][51] = 6;
        pixel_data[63][52] = 6;
        pixel_data[63][53] = 6;
        pixel_data[63][54] = 6;
        pixel_data[63][55] = 6;
        pixel_data[63][56] = 6;
        pixel_data[63][57] = 6;
        pixel_data[63][58] = 6;
        pixel_data[63][59] = 6;
        pixel_data[63][60] = 6;
        pixel_data[63][61] = 6;
        pixel_data[63][62] = 6;
        pixel_data[63][63] = 6;
        pixel_data[63][64] = 6;
        pixel_data[63][65] = 6;
        pixel_data[63][66] = 6;
        pixel_data[63][67] = 6;
        pixel_data[63][68] = 6;
        pixel_data[63][69] = 6;
        pixel_data[63][70] = 12;
        pixel_data[63][71] = 0;
        pixel_data[63][72] = 0;
        pixel_data[63][73] = 0;
        pixel_data[63][74] = 0;
        pixel_data[63][75] = 0;
        pixel_data[63][76] = 0;
        pixel_data[63][77] = 0;
        pixel_data[63][78] = 0;
        pixel_data[63][79] = 0;
        pixel_data[63][80] = 0;
        pixel_data[63][81] = 0;
        pixel_data[63][82] = 0;
        pixel_data[63][83] = 0;
        pixel_data[63][84] = 0;
        pixel_data[63][85] = 0;
        pixel_data[63][86] = 0;
        pixel_data[63][87] = 0;
        pixel_data[63][88] = 0;
        pixel_data[63][89] = 0;
        pixel_data[63][90] = 0;
        pixel_data[63][91] = 0;
        pixel_data[63][92] = 0;
        pixel_data[63][93] = 0;
        pixel_data[63][94] = 0;
        pixel_data[63][95] = 0;
        pixel_data[63][96] = 0;
        pixel_data[63][97] = 0;
        pixel_data[63][98] = 0;
        pixel_data[63][99] = 0; // y=63
        pixel_data[64][0] = 0;
        pixel_data[64][1] = 0;
        pixel_data[64][2] = 0;
        pixel_data[64][3] = 0;
        pixel_data[64][4] = 0;
        pixel_data[64][5] = 0;
        pixel_data[64][6] = 0;
        pixel_data[64][7] = 0;
        pixel_data[64][8] = 0;
        pixel_data[64][9] = 0;
        pixel_data[64][10] = 0;
        pixel_data[64][11] = 8;
        pixel_data[64][12] = 8;
        pixel_data[64][13] = 9;
        pixel_data[64][14] = 10;
        pixel_data[64][15] = 11;
        pixel_data[64][16] = 11;
        pixel_data[64][17] = 11;
        pixel_data[64][18] = 11;
        pixel_data[64][19] = 11;
        pixel_data[64][20] = 11;
        pixel_data[64][21] = 12;
        pixel_data[64][22] = 12;
        pixel_data[64][23] = 12;
        pixel_data[64][24] = 12;
        pixel_data[64][25] = 12;
        pixel_data[64][26] = 12;
        pixel_data[64][27] = 12;
        pixel_data[64][28] = 11;
        pixel_data[64][29] = 11;
        pixel_data[64][30] = 10;
        pixel_data[64][31] = 9;
        pixel_data[64][32] = 9;
        pixel_data[64][33] = 8;
        pixel_data[64][34] = 8;
        pixel_data[64][35] = 8;
        pixel_data[64][36] = 6;
        pixel_data[64][37] = 6;
        pixel_data[64][38] = 6;
        pixel_data[64][39] = 6;
        pixel_data[64][40] = 6;
        pixel_data[64][41] = 6;
        pixel_data[64][42] = 6;
        pixel_data[64][43] = 6;
        pixel_data[64][44] = 6;
        pixel_data[64][45] = 6;
        pixel_data[64][46] = 6;
        pixel_data[64][47] = 6;
        pixel_data[64][48] = 6;
        pixel_data[64][49] = 6;
        pixel_data[64][50] = 6;
        pixel_data[64][51] = 6;
        pixel_data[64][52] = 6;
        pixel_data[64][53] = 6;
        pixel_data[64][54] = 6;
        pixel_data[64][55] = 6;
        pixel_data[64][56] = 6;
        pixel_data[64][57] = 6;
        pixel_data[64][58] = 6;
        pixel_data[64][59] = 6;
        pixel_data[64][60] = 6;
        pixel_data[64][61] = 6;
        pixel_data[64][62] = 6;
        pixel_data[64][63] = 6;
        pixel_data[64][64] = 6;
        pixel_data[64][65] = 6;
        pixel_data[64][66] = 6;
        pixel_data[64][67] = 6;
        pixel_data[64][68] = 11;
        pixel_data[64][69] = 1;
        pixel_data[64][70] = 0;
        pixel_data[64][71] = 0;
        pixel_data[64][72] = 0;
        pixel_data[64][73] = 0;
        pixel_data[64][74] = 0;
        pixel_data[64][75] = 0;
        pixel_data[64][76] = 0;
        pixel_data[64][77] = 0;
        pixel_data[64][78] = 0;
        pixel_data[64][79] = 0;
        pixel_data[64][80] = 0;
        pixel_data[64][81] = 0;
        pixel_data[64][82] = 0;
        pixel_data[64][83] = 0;
        pixel_data[64][84] = 0;
        pixel_data[64][85] = 0;
        pixel_data[64][86] = 0;
        pixel_data[64][87] = 0;
        pixel_data[64][88] = 0;
        pixel_data[64][89] = 0;
        pixel_data[64][90] = 0;
        pixel_data[64][91] = 0;
        pixel_data[64][92] = 0;
        pixel_data[64][93] = 0;
        pixel_data[64][94] = 0;
        pixel_data[64][95] = 0;
        pixel_data[64][96] = 0;
        pixel_data[64][97] = 0;
        pixel_data[64][98] = 0;
        pixel_data[64][99] = 0; // y=64
        pixel_data[65][0] = 0;
        pixel_data[65][1] = 0;
        pixel_data[65][2] = 0;
        pixel_data[65][3] = 0;
        pixel_data[65][4] = 0;
        pixel_data[65][5] = 0;
        pixel_data[65][6] = 0;
        pixel_data[65][7] = 0;
        pixel_data[65][8] = 0;
        pixel_data[65][9] = 0;
        pixel_data[65][10] = 14;
        pixel_data[65][11] = 8;
        pixel_data[65][12] = 8;
        pixel_data[65][13] = 9;
        pixel_data[65][14] = 10;
        pixel_data[65][15] = 11;
        pixel_data[65][16] = 11;
        pixel_data[65][17] = 11;
        pixel_data[65][18] = 11;
        pixel_data[65][19] = 11;
        pixel_data[65][20] = 11;
        pixel_data[65][21] = 11;
        pixel_data[65][22] = 12;
        pixel_data[65][23] = 12;
        pixel_data[65][24] = 12;
        pixel_data[65][25] = 12;
        pixel_data[65][26] = 11;
        pixel_data[65][27] = 11;
        pixel_data[65][28] = 10;
        pixel_data[65][29] = 9;
        pixel_data[65][30] = 8;
        pixel_data[65][31] = 8;
        pixel_data[65][32] = 6;
        pixel_data[65][33] = 6;
        pixel_data[65][34] = 6;
        pixel_data[65][35] = 6;
        pixel_data[65][36] = 6;
        pixel_data[65][37] = 6;
        pixel_data[65][38] = 6;
        pixel_data[65][39] = 6;
        pixel_data[65][40] = 6;
        pixel_data[65][41] = 6;
        pixel_data[65][42] = 6;
        pixel_data[65][43] = 6;
        pixel_data[65][44] = 6;
        pixel_data[65][45] = 6;
        pixel_data[65][46] = 6;
        pixel_data[65][47] = 6;
        pixel_data[65][48] = 6;
        pixel_data[65][49] = 6;
        pixel_data[65][50] = 6;
        pixel_data[65][51] = 6;
        pixel_data[65][52] = 6;
        pixel_data[65][53] = 6;
        pixel_data[65][54] = 6;
        pixel_data[65][55] = 6;
        pixel_data[65][56] = 6;
        pixel_data[65][57] = 6;
        pixel_data[65][58] = 6;
        pixel_data[65][59] = 6;
        pixel_data[65][60] = 6;
        pixel_data[65][61] = 6;
        pixel_data[65][62] = 6;
        pixel_data[65][63] = 6;
        pixel_data[65][64] = 6;
        pixel_data[65][65] = 6;
        pixel_data[65][66] = 2;
        pixel_data[65][67] = 1;
        pixel_data[65][68] = 0;
        pixel_data[65][69] = 0;
        pixel_data[65][70] = 0;
        pixel_data[65][71] = 0;
        pixel_data[65][72] = 0;
        pixel_data[65][73] = 0;
        pixel_data[65][74] = 0;
        pixel_data[65][75] = 0;
        pixel_data[65][76] = 0;
        pixel_data[65][77] = 0;
        pixel_data[65][78] = 0;
        pixel_data[65][79] = 0;
        pixel_data[65][80] = 0;
        pixel_data[65][81] = 0;
        pixel_data[65][82] = 0;
        pixel_data[65][83] = 0;
        pixel_data[65][84] = 0;
        pixel_data[65][85] = 0;
        pixel_data[65][86] = 0;
        pixel_data[65][87] = 0;
        pixel_data[65][88] = 0;
        pixel_data[65][89] = 0;
        pixel_data[65][90] = 0;
        pixel_data[65][91] = 0;
        pixel_data[65][92] = 0;
        pixel_data[65][93] = 0;
        pixel_data[65][94] = 0;
        pixel_data[65][95] = 0;
        pixel_data[65][96] = 0;
        pixel_data[65][97] = 0;
        pixel_data[65][98] = 0;
        pixel_data[65][99] = 0; // y=65
        pixel_data[66][0] = 0;
        pixel_data[66][1] = 0;
        pixel_data[66][2] = 0;
        pixel_data[66][3] = 0;
        pixel_data[66][4] = 0;
        pixel_data[66][5] = 0;
        pixel_data[66][6] = 0;
        pixel_data[66][7] = 0;
        pixel_data[66][8] = 0;
        pixel_data[66][9] = 0;
        pixel_data[66][10] = 7;
        pixel_data[66][11] = 8;
        pixel_data[66][12] = 8;
        pixel_data[66][13] = 9;
        pixel_data[66][14] = 10;
        pixel_data[66][15] = 10;
        pixel_data[66][16] = 11;
        pixel_data[66][17] = 11;
        pixel_data[66][18] = 11;
        pixel_data[66][19] = 11;
        pixel_data[66][20] = 11;
        pixel_data[66][21] = 11;
        pixel_data[66][22] = 11;
        pixel_data[66][23] = 12;
        pixel_data[66][24] = 11;
        pixel_data[66][25] = 11;
        pixel_data[66][26] = 10;
        pixel_data[66][27] = 10;
        pixel_data[66][28] = 9;
        pixel_data[66][29] = 6;
        pixel_data[66][30] = 6;
        pixel_data[66][31] = 6;
        pixel_data[66][32] = 6;
        pixel_data[66][33] = 6;
        pixel_data[66][34] = 6;
        pixel_data[66][35] = 6;
        pixel_data[66][36] = 6;
        pixel_data[66][37] = 6;
        pixel_data[66][38] = 6;
        pixel_data[66][39] = 6;
        pixel_data[66][40] = 6;
        pixel_data[66][41] = 6;
        pixel_data[66][42] = 6;
        pixel_data[66][43] = 6;
        pixel_data[66][44] = 6;
        pixel_data[66][45] = 6;
        pixel_data[66][46] = 6;
        pixel_data[66][47] = 6;
        pixel_data[66][48] = 6;
        pixel_data[66][49] = 6;
        pixel_data[66][50] = 6;
        pixel_data[66][51] = 6;
        pixel_data[66][52] = 6;
        pixel_data[66][53] = 6;
        pixel_data[66][54] = 6;
        pixel_data[66][55] = 6;
        pixel_data[66][56] = 6;
        pixel_data[66][57] = 6;
        pixel_data[66][58] = 6;
        pixel_data[66][59] = 6;
        pixel_data[66][60] = 6;
        pixel_data[66][61] = 6;
        pixel_data[66][62] = 8;
        pixel_data[66][63] = 7;
        pixel_data[66][64] = 7;
        pixel_data[66][65] = 0;
        pixel_data[66][66] = 0;
        pixel_data[66][67] = 0;
        pixel_data[66][68] = 0;
        pixel_data[66][69] = 0;
        pixel_data[66][70] = 0;
        pixel_data[66][71] = 0;
        pixel_data[66][72] = 0;
        pixel_data[66][73] = 0;
        pixel_data[66][74] = 0;
        pixel_data[66][75] = 0;
        pixel_data[66][76] = 0;
        pixel_data[66][77] = 0;
        pixel_data[66][78] = 0;
        pixel_data[66][79] = 0;
        pixel_data[66][80] = 0;
        pixel_data[66][81] = 0;
        pixel_data[66][82] = 0;
        pixel_data[66][83] = 0;
        pixel_data[66][84] = 0;
        pixel_data[66][85] = 0;
        pixel_data[66][86] = 0;
        pixel_data[66][87] = 0;
        pixel_data[66][88] = 0;
        pixel_data[66][89] = 0;
        pixel_data[66][90] = 0;
        pixel_data[66][91] = 0;
        pixel_data[66][92] = 0;
        pixel_data[66][93] = 0;
        pixel_data[66][94] = 0;
        pixel_data[66][95] = 0;
        pixel_data[66][96] = 0;
        pixel_data[66][97] = 0;
        pixel_data[66][98] = 0;
        pixel_data[66][99] = 0; // y=66
        pixel_data[67][0] = 0;
        pixel_data[67][1] = 0;
        pixel_data[67][2] = 0;
        pixel_data[67][3] = 0;
        pixel_data[67][4] = 0;
        pixel_data[67][5] = 0;
        pixel_data[67][6] = 0;
        pixel_data[67][7] = 0;
        pixel_data[67][8] = 0;
        pixel_data[67][9] = 0;
        pixel_data[67][10] = 5;
        pixel_data[67][11] = 6;
        pixel_data[67][12] = 8;
        pixel_data[67][13] = 9;
        pixel_data[67][14] = 9;
        pixel_data[67][15] = 10;
        pixel_data[67][16] = 10;
        pixel_data[67][17] = 11;
        pixel_data[67][18] = 11;
        pixel_data[67][19] = 11;
        pixel_data[67][20] = 11;
        pixel_data[67][21] = 11;
        pixel_data[67][22] = 11;
        pixel_data[67][23] = 11;
        pixel_data[67][24] = 10;
        pixel_data[67][25] = 9;
        pixel_data[67][26] = 9;
        pixel_data[67][27] = 8;
        pixel_data[67][28] = 6;
        pixel_data[67][29] = 6;
        pixel_data[67][30] = 6;
        pixel_data[67][31] = 6;
        pixel_data[67][32] = 6;
        pixel_data[67][33] = 6;
        pixel_data[67][34] = 6;
        pixel_data[67][35] = 6;
        pixel_data[67][36] = 8;
        pixel_data[67][37] = 6;
        pixel_data[67][38] = 6;
        pixel_data[67][39] = 6;
        pixel_data[67][40] = 6;
        pixel_data[67][41] = 6;
        pixel_data[67][42] = 6;
        pixel_data[67][43] = 6;
        pixel_data[67][44] = 6;
        pixel_data[67][45] = 6;
        pixel_data[67][46] = 6;
        pixel_data[67][47] = 6;
        pixel_data[67][48] = 6;
        pixel_data[67][49] = 6;
        pixel_data[67][50] = 6;
        pixel_data[67][51] = 6;
        pixel_data[67][52] = 6;
        pixel_data[67][53] = 6;
        pixel_data[67][54] = 8;
        pixel_data[67][55] = 8;
        pixel_data[67][56] = 5;
        pixel_data[67][57] = 5;
        pixel_data[67][58] = 2;
        pixel_data[67][59] = 2;
        pixel_data[67][60] = 15;
        pixel_data[67][61] = 0;
        pixel_data[67][62] = 0;
        pixel_data[67][63] = 0;
        pixel_data[67][64] = 0;
        pixel_data[67][65] = 0;
        pixel_data[67][66] = 0;
        pixel_data[67][67] = 0;
        pixel_data[67][68] = 0;
        pixel_data[67][69] = 0;
        pixel_data[67][70] = 0;
        pixel_data[67][71] = 0;
        pixel_data[67][72] = 0;
        pixel_data[67][73] = 0;
        pixel_data[67][74] = 0;
        pixel_data[67][75] = 0;
        pixel_data[67][76] = 0;
        pixel_data[67][77] = 0;
        pixel_data[67][78] = 0;
        pixel_data[67][79] = 0;
        pixel_data[67][80] = 0;
        pixel_data[67][81] = 0;
        pixel_data[67][82] = 0;
        pixel_data[67][83] = 0;
        pixel_data[67][84] = 0;
        pixel_data[67][85] = 0;
        pixel_data[67][86] = 0;
        pixel_data[67][87] = 0;
        pixel_data[67][88] = 0;
        pixel_data[67][89] = 0;
        pixel_data[67][90] = 0;
        pixel_data[67][91] = 0;
        pixel_data[67][92] = 0;
        pixel_data[67][93] = 0;
        pixel_data[67][94] = 0;
        pixel_data[67][95] = 0;
        pixel_data[67][96] = 0;
        pixel_data[67][97] = 0;
        pixel_data[67][98] = 0;
        pixel_data[67][99] = 0; // y=67
        pixel_data[68][0] = 0;
        pixel_data[68][1] = 0;
        pixel_data[68][2] = 0;
        pixel_data[68][3] = 0;
        pixel_data[68][4] = 0;
        pixel_data[68][5] = 0;
        pixel_data[68][6] = 0;
        pixel_data[68][7] = 0;
        pixel_data[68][8] = 0;
        pixel_data[68][9] = 15;
        pixel_data[68][10] = 6;
        pixel_data[68][11] = 6;
        pixel_data[68][12] = 6;
        pixel_data[68][13] = 8;
        pixel_data[68][14] = 9;
        pixel_data[68][15] = 9;
        pixel_data[68][16] = 10;
        pixel_data[68][17] = 10;
        pixel_data[68][18] = 11;
        pixel_data[68][19] = 11;
        pixel_data[68][20] = 11;
        pixel_data[68][21] = 11;
        pixel_data[68][22] = 11;
        pixel_data[68][23] = 10;
        pixel_data[68][24] = 9;
        pixel_data[68][25] = 8;
        pixel_data[68][26] = 6;
        pixel_data[68][27] = 6;
        pixel_data[68][28] = 6;
        pixel_data[68][29] = 6;
        pixel_data[68][30] = 6;
        pixel_data[68][31] = 6;
        pixel_data[68][32] = 6;
        pixel_data[68][33] = 5;
        pixel_data[68][34] = 2;
        pixel_data[68][35] = 5;
        pixel_data[68][36] = 2;
        pixel_data[68][37] = 14;
        pixel_data[68][38] = 7;
        pixel_data[68][39] = 7;
        pixel_data[68][40] = 7;
        pixel_data[68][41] = 12;
        pixel_data[68][42] = 7;
        pixel_data[68][43] = 7;
        pixel_data[68][44] = 7;
        pixel_data[68][45] = 12;
        pixel_data[68][46] = 7;
        pixel_data[68][47] = 14;
        pixel_data[68][48] = 15;
        pixel_data[68][49] = 1;
        pixel_data[68][50] = 0;
        pixel_data[68][51] = 0;
        pixel_data[68][52] = 1;
        pixel_data[68][53] = 0;
        pixel_data[68][54] = 0;
        pixel_data[68][55] = 0;
        pixel_data[68][56] = 0;
        pixel_data[68][57] = 0;
        pixel_data[68][58] = 0;
        pixel_data[68][59] = 0;
        pixel_data[68][60] = 0;
        pixel_data[68][61] = 0;
        pixel_data[68][62] = 0;
        pixel_data[68][63] = 0;
        pixel_data[68][64] = 0;
        pixel_data[68][65] = 0;
        pixel_data[68][66] = 0;
        pixel_data[68][67] = 0;
        pixel_data[68][68] = 0;
        pixel_data[68][69] = 0;
        pixel_data[68][70] = 0;
        pixel_data[68][71] = 0;
        pixel_data[68][72] = 0;
        pixel_data[68][73] = 0;
        pixel_data[68][74] = 0;
        pixel_data[68][75] = 0;
        pixel_data[68][76] = 0;
        pixel_data[68][77] = 0;
        pixel_data[68][78] = 0;
        pixel_data[68][79] = 0;
        pixel_data[68][80] = 0;
        pixel_data[68][81] = 0;
        pixel_data[68][82] = 0;
        pixel_data[68][83] = 0;
        pixel_data[68][84] = 0;
        pixel_data[68][85] = 0;
        pixel_data[68][86] = 0;
        pixel_data[68][87] = 0;
        pixel_data[68][88] = 0;
        pixel_data[68][89] = 0;
        pixel_data[68][90] = 0;
        pixel_data[68][91] = 0;
        pixel_data[68][92] = 0;
        pixel_data[68][93] = 0;
        pixel_data[68][94] = 0;
        pixel_data[68][95] = 0;
        pixel_data[68][96] = 0;
        pixel_data[68][97] = 0;
        pixel_data[68][98] = 0;
        pixel_data[68][99] = 0; // y=68
        pixel_data[69][0] = 0;
        pixel_data[69][1] = 0;
        pixel_data[69][2] = 0;
        pixel_data[69][3] = 0;
        pixel_data[69][4] = 0;
        pixel_data[69][5] = 0;
        pixel_data[69][6] = 0;
        pixel_data[69][7] = 0;
        pixel_data[69][8] = 0;
        pixel_data[69][9] = 4;
        pixel_data[69][10] = 6;
        pixel_data[69][11] = 6;
        pixel_data[69][12] = 6;
        pixel_data[69][13] = 6;
        pixel_data[69][14] = 8;
        pixel_data[69][15] = 9;
        pixel_data[69][16] = 9;
        pixel_data[69][17] = 10;
        pixel_data[69][18] = 10;
        pixel_data[69][19] = 10;
        pixel_data[69][20] = 10;
        pixel_data[69][21] = 10;
        pixel_data[69][22] = 9;
        pixel_data[69][23] = 9;
        pixel_data[69][24] = 8;
        pixel_data[69][25] = 6;
        pixel_data[69][26] = 6;
        pixel_data[69][27] = 6;
        pixel_data[69][28] = 6;
        pixel_data[69][29] = 8;
        pixel_data[69][30] = 7;
        pixel_data[69][31] = 7;
        pixel_data[69][32] = 0;
        pixel_data[69][33] = 0;
        pixel_data[69][34] = 0;
        pixel_data[69][35] = 0;
        pixel_data[69][36] = 0;
        pixel_data[69][37] = 0;
        pixel_data[69][38] = 0;
        pixel_data[69][39] = 0;
        pixel_data[69][40] = 0;
        pixel_data[69][41] = 0;
        pixel_data[69][42] = 0;
        pixel_data[69][43] = 0;
        pixel_data[69][44] = 0;
        pixel_data[69][45] = 0;
        pixel_data[69][46] = 0;
        pixel_data[69][47] = 0;
        pixel_data[69][48] = 0;
        pixel_data[69][49] = 0;
        pixel_data[69][50] = 0;
        pixel_data[69][51] = 0;
        pixel_data[69][52] = 0;
        pixel_data[69][53] = 0;
        pixel_data[69][54] = 0;
        pixel_data[69][55] = 0;
        pixel_data[69][56] = 0;
        pixel_data[69][57] = 0;
        pixel_data[69][58] = 0;
        pixel_data[69][59] = 0;
        pixel_data[69][60] = 0;
        pixel_data[69][61] = 0;
        pixel_data[69][62] = 0;
        pixel_data[69][63] = 0;
        pixel_data[69][64] = 0;
        pixel_data[69][65] = 0;
        pixel_data[69][66] = 0;
        pixel_data[69][67] = 0;
        pixel_data[69][68] = 0;
        pixel_data[69][69] = 0;
        pixel_data[69][70] = 0;
        pixel_data[69][71] = 0;
        pixel_data[69][72] = 0;
        pixel_data[69][73] = 0;
        pixel_data[69][74] = 0;
        pixel_data[69][75] = 0;
        pixel_data[69][76] = 0;
        pixel_data[69][77] = 0;
        pixel_data[69][78] = 0;
        pixel_data[69][79] = 0;
        pixel_data[69][80] = 0;
        pixel_data[69][81] = 0;
        pixel_data[69][82] = 0;
        pixel_data[69][83] = 0;
        pixel_data[69][84] = 0;
        pixel_data[69][85] = 0;
        pixel_data[69][86] = 0;
        pixel_data[69][87] = 0;
        pixel_data[69][88] = 0;
        pixel_data[69][89] = 0;
        pixel_data[69][90] = 0;
        pixel_data[69][91] = 0;
        pixel_data[69][92] = 0;
        pixel_data[69][93] = 0;
        pixel_data[69][94] = 0;
        pixel_data[69][95] = 0;
        pixel_data[69][96] = 0;
        pixel_data[69][97] = 0;
        pixel_data[69][98] = 0;
        pixel_data[69][99] = 0; // y=69
        pixel_data[70][0] = 0;
        pixel_data[70][1] = 0;
        pixel_data[70][2] = 0;
        pixel_data[70][3] = 0;
        pixel_data[70][4] = 0;
        pixel_data[70][5] = 0;
        pixel_data[70][6] = 0;
        pixel_data[70][7] = 0;
        pixel_data[70][8] = 0;
        pixel_data[70][9] = 8;
        pixel_data[70][10] = 6;
        pixel_data[70][11] = 6;
        pixel_data[70][12] = 6;
        pixel_data[70][13] = 6;
        pixel_data[70][14] = 6;
        pixel_data[70][15] = 8;
        pixel_data[70][16] = 8;
        pixel_data[70][17] = 9;
        pixel_data[70][18] = 9;
        pixel_data[70][19] = 9;
        pixel_data[70][20] = 9;
        pixel_data[70][21] = 9;
        pixel_data[70][22] = 8;
        pixel_data[70][23] = 6;
        pixel_data[70][24] = 6;
        pixel_data[70][25] = 6;
        pixel_data[70][26] = 6;
        pixel_data[70][27] = 6;
        pixel_data[70][28] = 5;
        pixel_data[70][29] = 7;
        pixel_data[70][30] = 0;
        pixel_data[70][31] = 0;
        pixel_data[70][32] = 0;
        pixel_data[70][33] = 0;
        pixel_data[70][34] = 0;
        pixel_data[70][35] = 0;
        pixel_data[70][36] = 0;
        pixel_data[70][37] = 0;
        pixel_data[70][38] = 0;
        pixel_data[70][39] = 0;
        pixel_data[70][40] = 0;
        pixel_data[70][41] = 0;
        pixel_data[70][42] = 0;
        pixel_data[70][43] = 0;
        pixel_data[70][44] = 0;
        pixel_data[70][45] = 0;
        pixel_data[70][46] = 0;
        pixel_data[70][47] = 0;
        pixel_data[70][48] = 0;
        pixel_data[70][49] = 0;
        pixel_data[70][50] = 0;
        pixel_data[70][51] = 0;
        pixel_data[70][52] = 0;
        pixel_data[70][53] = 0;
        pixel_data[70][54] = 0;
        pixel_data[70][55] = 0;
        pixel_data[70][56] = 0;
        pixel_data[70][57] = 0;
        pixel_data[70][58] = 0;
        pixel_data[70][59] = 0;
        pixel_data[70][60] = 0;
        pixel_data[70][61] = 0;
        pixel_data[70][62] = 0;
        pixel_data[70][63] = 0;
        pixel_data[70][64] = 0;
        pixel_data[70][65] = 0;
        pixel_data[70][66] = 0;
        pixel_data[70][67] = 0;
        pixel_data[70][68] = 0;
        pixel_data[70][69] = 0;
        pixel_data[70][70] = 0;
        pixel_data[70][71] = 0;
        pixel_data[70][72] = 0;
        pixel_data[70][73] = 0;
        pixel_data[70][74] = 0;
        pixel_data[70][75] = 0;
        pixel_data[70][76] = 0;
        pixel_data[70][77] = 0;
        pixel_data[70][78] = 0;
        pixel_data[70][79] = 0;
        pixel_data[70][80] = 0;
        pixel_data[70][81] = 0;
        pixel_data[70][82] = 0;
        pixel_data[70][83] = 0;
        pixel_data[70][84] = 0;
        pixel_data[70][85] = 0;
        pixel_data[70][86] = 0;
        pixel_data[70][87] = 0;
        pixel_data[70][88] = 0;
        pixel_data[70][89] = 0;
        pixel_data[70][90] = 0;
        pixel_data[70][91] = 0;
        pixel_data[70][92] = 0;
        pixel_data[70][93] = 0;
        pixel_data[70][94] = 0;
        pixel_data[70][95] = 0;
        pixel_data[70][96] = 0;
        pixel_data[70][97] = 0;
        pixel_data[70][98] = 0;
        pixel_data[70][99] = 0; // y=70
        pixel_data[71][0] = 0;
        pixel_data[71][1] = 0;
        pixel_data[71][2] = 0;
        pixel_data[71][3] = 0;
        pixel_data[71][4] = 0;
        pixel_data[71][5] = 0;
        pixel_data[71][6] = 0;
        pixel_data[71][7] = 0;
        pixel_data[71][8] = 7;
        pixel_data[71][9] = 6;
        pixel_data[71][10] = 6;
        pixel_data[71][11] = 6;
        pixel_data[71][12] = 6;
        pixel_data[71][13] = 6;
        pixel_data[71][14] = 6;
        pixel_data[71][15] = 6;
        pixel_data[71][16] = 6;
        pixel_data[71][17] = 8;
        pixel_data[71][18] = 8;
        pixel_data[71][19] = 8;
        pixel_data[71][20] = 8;
        pixel_data[71][21] = 8;
        pixel_data[71][22] = 6;
        pixel_data[71][23] = 6;
        pixel_data[71][24] = 6;
        pixel_data[71][25] = 6;
        pixel_data[71][26] = 6;
        pixel_data[71][27] = 7;
        pixel_data[71][28] = 0;
        pixel_data[71][29] = 0;
        pixel_data[71][30] = 0;
        pixel_data[71][31] = 0;
        pixel_data[71][32] = 0;
        pixel_data[71][33] = 0;
        pixel_data[71][34] = 0;
        pixel_data[71][35] = 0;
        pixel_data[71][36] = 0;
        pixel_data[71][37] = 0;
        pixel_data[71][38] = 0;
        pixel_data[71][39] = 0;
        pixel_data[71][40] = 0;
        pixel_data[71][41] = 0;
        pixel_data[71][42] = 0;
        pixel_data[71][43] = 0;
        pixel_data[71][44] = 0;
        pixel_data[71][45] = 0;
        pixel_data[71][46] = 0;
        pixel_data[71][47] = 0;
        pixel_data[71][48] = 0;
        pixel_data[71][49] = 0;
        pixel_data[71][50] = 0;
        pixel_data[71][51] = 0;
        pixel_data[71][52] = 0;
        pixel_data[71][53] = 0;
        pixel_data[71][54] = 0;
        pixel_data[71][55] = 0;
        pixel_data[71][56] = 0;
        pixel_data[71][57] = 0;
        pixel_data[71][58] = 0;
        pixel_data[71][59] = 0;
        pixel_data[71][60] = 0;
        pixel_data[71][61] = 0;
        pixel_data[71][62] = 0;
        pixel_data[71][63] = 0;
        pixel_data[71][64] = 0;
        pixel_data[71][65] = 0;
        pixel_data[71][66] = 0;
        pixel_data[71][67] = 0;
        pixel_data[71][68] = 0;
        pixel_data[71][69] = 0;
        pixel_data[71][70] = 0;
        pixel_data[71][71] = 0;
        pixel_data[71][72] = 0;
        pixel_data[71][73] = 0;
        pixel_data[71][74] = 0;
        pixel_data[71][75] = 0;
        pixel_data[71][76] = 0;
        pixel_data[71][77] = 0;
        pixel_data[71][78] = 0;
        pixel_data[71][79] = 0;
        pixel_data[71][80] = 0;
        pixel_data[71][81] = 0;
        pixel_data[71][82] = 0;
        pixel_data[71][83] = 0;
        pixel_data[71][84] = 0;
        pixel_data[71][85] = 0;
        pixel_data[71][86] = 0;
        pixel_data[71][87] = 0;
        pixel_data[71][88] = 0;
        pixel_data[71][89] = 0;
        pixel_data[71][90] = 0;
        pixel_data[71][91] = 0;
        pixel_data[71][92] = 0;
        pixel_data[71][93] = 0;
        pixel_data[71][94] = 0;
        pixel_data[71][95] = 0;
        pixel_data[71][96] = 0;
        pixel_data[71][97] = 0;
        pixel_data[71][98] = 0;
        pixel_data[71][99] = 0; // y=71
        pixel_data[72][0] = 0;
        pixel_data[72][1] = 0;
        pixel_data[72][2] = 0;
        pixel_data[72][3] = 0;
        pixel_data[72][4] = 0;
        pixel_data[72][5] = 0;
        pixel_data[72][6] = 0;
        pixel_data[72][7] = 0;
        pixel_data[72][8] = 2;
        pixel_data[72][9] = 6;
        pixel_data[72][10] = 6;
        pixel_data[72][11] = 6;
        pixel_data[72][12] = 6;
        pixel_data[72][13] = 6;
        pixel_data[72][14] = 6;
        pixel_data[72][15] = 6;
        pixel_data[72][16] = 6;
        pixel_data[72][17] = 6;
        pixel_data[72][18] = 6;
        pixel_data[72][19] = 6;
        pixel_data[72][20] = 6;
        pixel_data[72][21] = 6;
        pixel_data[72][22] = 6;
        pixel_data[72][23] = 6;
        pixel_data[72][24] = 6;
        pixel_data[72][25] = 2;
        pixel_data[72][26] = 0;
        pixel_data[72][27] = 0;
        pixel_data[72][28] = 0;
        pixel_data[72][29] = 0;
        pixel_data[72][30] = 0;
        pixel_data[72][31] = 0;
        pixel_data[72][32] = 0;
        pixel_data[72][33] = 0;
        pixel_data[72][34] = 0;
        pixel_data[72][35] = 0;
        pixel_data[72][36] = 0;
        pixel_data[72][37] = 0;
        pixel_data[72][38] = 0;
        pixel_data[72][39] = 0;
        pixel_data[72][40] = 0;
        pixel_data[72][41] = 0;
        pixel_data[72][42] = 0;
        pixel_data[72][43] = 0;
        pixel_data[72][44] = 0;
        pixel_data[72][45] = 0;
        pixel_data[72][46] = 0;
        pixel_data[72][47] = 0;
        pixel_data[72][48] = 0;
        pixel_data[72][49] = 0;
        pixel_data[72][50] = 0;
        pixel_data[72][51] = 0;
        pixel_data[72][52] = 0;
        pixel_data[72][53] = 0;
        pixel_data[72][54] = 0;
        pixel_data[72][55] = 0;
        pixel_data[72][56] = 0;
        pixel_data[72][57] = 0;
        pixel_data[72][58] = 0;
        pixel_data[72][59] = 0;
        pixel_data[72][60] = 0;
        pixel_data[72][61] = 0;
        pixel_data[72][62] = 0;
        pixel_data[72][63] = 0;
        pixel_data[72][64] = 0;
        pixel_data[72][65] = 0;
        pixel_data[72][66] = 0;
        pixel_data[72][67] = 0;
        pixel_data[72][68] = 0;
        pixel_data[72][69] = 0;
        pixel_data[72][70] = 0;
        pixel_data[72][71] = 0;
        pixel_data[72][72] = 0;
        pixel_data[72][73] = 0;
        pixel_data[72][74] = 0;
        pixel_data[72][75] = 0;
        pixel_data[72][76] = 0;
        pixel_data[72][77] = 0;
        pixel_data[72][78] = 0;
        pixel_data[72][79] = 0;
        pixel_data[72][80] = 0;
        pixel_data[72][81] = 0;
        pixel_data[72][82] = 0;
        pixel_data[72][83] = 0;
        pixel_data[72][84] = 0;
        pixel_data[72][85] = 0;
        pixel_data[72][86] = 0;
        pixel_data[72][87] = 0;
        pixel_data[72][88] = 0;
        pixel_data[72][89] = 0;
        pixel_data[72][90] = 0;
        pixel_data[72][91] = 0;
        pixel_data[72][92] = 0;
        pixel_data[72][93] = 0;
        pixel_data[72][94] = 0;
        pixel_data[72][95] = 0;
        pixel_data[72][96] = 0;
        pixel_data[72][97] = 0;
        pixel_data[72][98] = 0;
        pixel_data[72][99] = 0; // y=72
        pixel_data[73][0] = 0;
        pixel_data[73][1] = 0;
        pixel_data[73][2] = 0;
        pixel_data[73][3] = 0;
        pixel_data[73][4] = 0;
        pixel_data[73][5] = 0;
        pixel_data[73][6] = 0;
        pixel_data[73][7] = 0;
        pixel_data[73][8] = 2;
        pixel_data[73][9] = 8;
        pixel_data[73][10] = 6;
        pixel_data[73][11] = 6;
        pixel_data[73][12] = 6;
        pixel_data[73][13] = 6;
        pixel_data[73][14] = 6;
        pixel_data[73][15] = 6;
        pixel_data[73][16] = 6;
        pixel_data[73][17] = 6;
        pixel_data[73][18] = 6;
        pixel_data[73][19] = 6;
        pixel_data[73][20] = 6;
        pixel_data[73][21] = 6;
        pixel_data[73][22] = 8;
        pixel_data[73][23] = 11;
        pixel_data[73][24] = 0;
        pixel_data[73][25] = 0;
        pixel_data[73][26] = 0;
        pixel_data[73][27] = 0;
        pixel_data[73][28] = 0;
        pixel_data[73][29] = 0;
        pixel_data[73][30] = 0;
        pixel_data[73][31] = 0;
        pixel_data[73][32] = 0;
        pixel_data[73][33] = 0;
        pixel_data[73][34] = 0;
        pixel_data[73][35] = 0;
        pixel_data[73][36] = 0;
        pixel_data[73][37] = 0;
        pixel_data[73][38] = 0;
        pixel_data[73][39] = 0;
        pixel_data[73][40] = 0;
        pixel_data[73][41] = 0;
        pixel_data[73][42] = 0;
        pixel_data[73][43] = 0;
        pixel_data[73][44] = 0;
        pixel_data[73][45] = 0;
        pixel_data[73][46] = 0;
        pixel_data[73][47] = 0;
        pixel_data[73][48] = 0;
        pixel_data[73][49] = 0;
        pixel_data[73][50] = 0;
        pixel_data[73][51] = 0;
        pixel_data[73][52] = 0;
        pixel_data[73][53] = 0;
        pixel_data[73][54] = 0;
        pixel_data[73][55] = 0;
        pixel_data[73][56] = 0;
        pixel_data[73][57] = 0;
        pixel_data[73][58] = 0;
        pixel_data[73][59] = 0;
        pixel_data[73][60] = 0;
        pixel_data[73][61] = 0;
        pixel_data[73][62] = 0;
        pixel_data[73][63] = 0;
        pixel_data[73][64] = 0;
        pixel_data[73][65] = 0;
        pixel_data[73][66] = 0;
        pixel_data[73][67] = 0;
        pixel_data[73][68] = 0;
        pixel_data[73][69] = 0;
        pixel_data[73][70] = 0;
        pixel_data[73][71] = 0;
        pixel_data[73][72] = 0;
        pixel_data[73][73] = 0;
        pixel_data[73][74] = 0;
        pixel_data[73][75] = 0;
        pixel_data[73][76] = 0;
        pixel_data[73][77] = 0;
        pixel_data[73][78] = 0;
        pixel_data[73][79] = 0;
        pixel_data[73][80] = 0;
        pixel_data[73][81] = 0;
        pixel_data[73][82] = 0;
        pixel_data[73][83] = 0;
        pixel_data[73][84] = 0;
        pixel_data[73][85] = 0;
        pixel_data[73][86] = 0;
        pixel_data[73][87] = 0;
        pixel_data[73][88] = 0;
        pixel_data[73][89] = 0;
        pixel_data[73][90] = 0;
        pixel_data[73][91] = 0;
        pixel_data[73][92] = 0;
        pixel_data[73][93] = 0;
        pixel_data[73][94] = 0;
        pixel_data[73][95] = 0;
        pixel_data[73][96] = 0;
        pixel_data[73][97] = 0;
        pixel_data[73][98] = 0;
        pixel_data[73][99] = 0; // y=73
        pixel_data[74][0] = 0;
        pixel_data[74][1] = 0;
        pixel_data[74][2] = 0;
        pixel_data[74][3] = 0;
        pixel_data[74][4] = 0;
        pixel_data[74][5] = 0;
        pixel_data[74][6] = 0;
        pixel_data[74][7] = 0;
        pixel_data[74][8] = 7;
        pixel_data[74][9] = 6;
        pixel_data[74][10] = 6;
        pixel_data[74][11] = 6;
        pixel_data[74][12] = 6;
        pixel_data[74][13] = 6;
        pixel_data[74][14] = 6;
        pixel_data[74][15] = 6;
        pixel_data[74][16] = 6;
        pixel_data[74][17] = 6;
        pixel_data[74][18] = 6;
        pixel_data[74][19] = 6;
        pixel_data[74][20] = 6;
        pixel_data[74][21] = 8;
        pixel_data[74][22] = 0;
        pixel_data[74][23] = 0;
        pixel_data[74][24] = 0;
        pixel_data[74][25] = 0;
        pixel_data[74][26] = 0;
        pixel_data[74][27] = 0;
        pixel_data[74][28] = 0;
        pixel_data[74][29] = 0;
        pixel_data[74][30] = 0;
        pixel_data[74][31] = 0;
        pixel_data[74][32] = 0;
        pixel_data[74][33] = 0;
        pixel_data[74][34] = 0;
        pixel_data[74][35] = 0;
        pixel_data[74][36] = 0;
        pixel_data[74][37] = 0;
        pixel_data[74][38] = 0;
        pixel_data[74][39] = 0;
        pixel_data[74][40] = 0;
        pixel_data[74][41] = 0;
        pixel_data[74][42] = 0;
        pixel_data[74][43] = 0;
        pixel_data[74][44] = 0;
        pixel_data[74][45] = 0;
        pixel_data[74][46] = 0;
        pixel_data[74][47] = 0;
        pixel_data[74][48] = 0;
        pixel_data[74][49] = 0;
        pixel_data[74][50] = 0;
        pixel_data[74][51] = 0;
        pixel_data[74][52] = 0;
        pixel_data[74][53] = 0;
        pixel_data[74][54] = 0;
        pixel_data[74][55] = 0;
        pixel_data[74][56] = 0;
        pixel_data[74][57] = 0;
        pixel_data[74][58] = 0;
        pixel_data[74][59] = 0;
        pixel_data[74][60] = 0;
        pixel_data[74][61] = 0;
        pixel_data[74][62] = 0;
        pixel_data[74][63] = 0;
        pixel_data[74][64] = 0;
        pixel_data[74][65] = 0;
        pixel_data[74][66] = 0;
        pixel_data[74][67] = 0;
        pixel_data[74][68] = 0;
        pixel_data[74][69] = 0;
        pixel_data[74][70] = 0;
        pixel_data[74][71] = 0;
        pixel_data[74][72] = 0;
        pixel_data[74][73] = 0;
        pixel_data[74][74] = 0;
        pixel_data[74][75] = 0;
        pixel_data[74][76] = 0;
        pixel_data[74][77] = 0;
        pixel_data[74][78] = 0;
        pixel_data[74][79] = 0;
        pixel_data[74][80] = 0;
        pixel_data[74][81] = 0;
        pixel_data[74][82] = 0;
        pixel_data[74][83] = 0;
        pixel_data[74][84] = 0;
        pixel_data[74][85] = 0;
        pixel_data[74][86] = 0;
        pixel_data[74][87] = 0;
        pixel_data[74][88] = 0;
        pixel_data[74][89] = 0;
        pixel_data[74][90] = 0;
        pixel_data[74][91] = 0;
        pixel_data[74][92] = 0;
        pixel_data[74][93] = 0;
        pixel_data[74][94] = 0;
        pixel_data[74][95] = 0;
        pixel_data[74][96] = 0;
        pixel_data[74][97] = 0;
        pixel_data[74][98] = 0;
        pixel_data[74][99] = 0; // y=74
        pixel_data[75][0] = 0;
        pixel_data[75][1] = 0;
        pixel_data[75][2] = 0;
        pixel_data[75][3] = 0;
        pixel_data[75][4] = 0;
        pixel_data[75][5] = 0;
        pixel_data[75][6] = 0;
        pixel_data[75][7] = 0;
        pixel_data[75][8] = 0;
        pixel_data[75][9] = 12;
        pixel_data[75][10] = 6;
        pixel_data[75][11] = 6;
        pixel_data[75][12] = 6;
        pixel_data[75][13] = 6;
        pixel_data[75][14] = 6;
        pixel_data[75][15] = 6;
        pixel_data[75][16] = 6;
        pixel_data[75][17] = 6;
        pixel_data[75][18] = 6;
        pixel_data[75][19] = 6;
        pixel_data[75][20] = 8;
        pixel_data[75][21] = 0;
        pixel_data[75][22] = 0;
        pixel_data[75][23] = 0;
        pixel_data[75][24] = 0;
        pixel_data[75][25] = 0;
        pixel_data[75][26] = 0;
        pixel_data[75][27] = 0;
        pixel_data[75][28] = 0;
        pixel_data[75][29] = 0;
        pixel_data[75][30] = 0;
        pixel_data[75][31] = 0;
        pixel_data[75][32] = 0;
        pixel_data[75][33] = 0;
        pixel_data[75][34] = 0;
        pixel_data[75][35] = 0;
        pixel_data[75][36] = 0;
        pixel_data[75][37] = 0;
        pixel_data[75][38] = 0;
        pixel_data[75][39] = 0;
        pixel_data[75][40] = 0;
        pixel_data[75][41] = 0;
        pixel_data[75][42] = 0;
        pixel_data[75][43] = 0;
        pixel_data[75][44] = 0;
        pixel_data[75][45] = 0;
        pixel_data[75][46] = 0;
        pixel_data[75][47] = 0;
        pixel_data[75][48] = 0;
        pixel_data[75][49] = 0;
        pixel_data[75][50] = 0;
        pixel_data[75][51] = 0;
        pixel_data[75][52] = 0;
        pixel_data[75][53] = 0;
        pixel_data[75][54] = 0;
        pixel_data[75][55] = 0;
        pixel_data[75][56] = 0;
        pixel_data[75][57] = 0;
        pixel_data[75][58] = 0;
        pixel_data[75][59] = 0;
        pixel_data[75][60] = 0;
        pixel_data[75][61] = 0;
        pixel_data[75][62] = 0;
        pixel_data[75][63] = 0;
        pixel_data[75][64] = 0;
        pixel_data[75][65] = 0;
        pixel_data[75][66] = 0;
        pixel_data[75][67] = 0;
        pixel_data[75][68] = 0;
        pixel_data[75][69] = 0;
        pixel_data[75][70] = 0;
        pixel_data[75][71] = 0;
        pixel_data[75][72] = 0;
        pixel_data[75][73] = 0;
        pixel_data[75][74] = 0;
        pixel_data[75][75] = 0;
        pixel_data[75][76] = 0;
        pixel_data[75][77] = 0;
        pixel_data[75][78] = 0;
        pixel_data[75][79] = 0;
        pixel_data[75][80] = 0;
        pixel_data[75][81] = 0;
        pixel_data[75][82] = 0;
        pixel_data[75][83] = 0;
        pixel_data[75][84] = 0;
        pixel_data[75][85] = 0;
        pixel_data[75][86] = 0;
        pixel_data[75][87] = 0;
        pixel_data[75][88] = 0;
        pixel_data[75][89] = 0;
        pixel_data[75][90] = 0;
        pixel_data[75][91] = 0;
        pixel_data[75][92] = 0;
        pixel_data[75][93] = 0;
        pixel_data[75][94] = 0;
        pixel_data[75][95] = 0;
        pixel_data[75][96] = 0;
        pixel_data[75][97] = 0;
        pixel_data[75][98] = 0;
        pixel_data[75][99] = 0; // y=75
        pixel_data[76][0] = 0;
        pixel_data[76][1] = 0;
        pixel_data[76][2] = 0;
        pixel_data[76][3] = 0;
        pixel_data[76][4] = 0;
        pixel_data[76][5] = 0;
        pixel_data[76][6] = 0;
        pixel_data[76][7] = 0;
        pixel_data[76][8] = 0;
        pixel_data[76][9] = 0;
        pixel_data[76][10] = 11;
        pixel_data[76][11] = 6;
        pixel_data[76][12] = 6;
        pixel_data[76][13] = 6;
        pixel_data[76][14] = 6;
        pixel_data[76][15] = 6;
        pixel_data[76][16] = 6;
        pixel_data[76][17] = 6;
        pixel_data[76][18] = 8;
        pixel_data[76][19] = 6;
        pixel_data[76][20] = 0;
        pixel_data[76][21] = 0;
        pixel_data[76][22] = 0;
        pixel_data[76][23] = 0;
        pixel_data[76][24] = 0;
        pixel_data[76][25] = 0;
        pixel_data[76][26] = 0;
        pixel_data[76][27] = 0;
        pixel_data[76][28] = 0;
        pixel_data[76][29] = 0;
        pixel_data[76][30] = 0;
        pixel_data[76][31] = 0;
        pixel_data[76][32] = 0;
        pixel_data[76][33] = 0;
        pixel_data[76][34] = 0;
        pixel_data[76][35] = 0;
        pixel_data[76][36] = 0;
        pixel_data[76][37] = 0;
        pixel_data[76][38] = 0;
        pixel_data[76][39] = 0;
        pixel_data[76][40] = 0;
        pixel_data[76][41] = 0;
        pixel_data[76][42] = 0;
        pixel_data[76][43] = 0;
        pixel_data[76][44] = 0;
        pixel_data[76][45] = 0;
        pixel_data[76][46] = 0;
        pixel_data[76][47] = 0;
        pixel_data[76][48] = 0;
        pixel_data[76][49] = 0;
        pixel_data[76][50] = 0;
        pixel_data[76][51] = 0;
        pixel_data[76][52] = 0;
        pixel_data[76][53] = 0;
        pixel_data[76][54] = 0;
        pixel_data[76][55] = 0;
        pixel_data[76][56] = 0;
        pixel_data[76][57] = 0;
        pixel_data[76][58] = 0;
        pixel_data[76][59] = 0;
        pixel_data[76][60] = 0;
        pixel_data[76][61] = 0;
        pixel_data[76][62] = 0;
        pixel_data[76][63] = 0;
        pixel_data[76][64] = 0;
        pixel_data[76][65] = 0;
        pixel_data[76][66] = 0;
        pixel_data[76][67] = 0;
        pixel_data[76][68] = 0;
        pixel_data[76][69] = 0;
        pixel_data[76][70] = 0;
        pixel_data[76][71] = 0;
        pixel_data[76][72] = 0;
        pixel_data[76][73] = 0;
        pixel_data[76][74] = 0;
        pixel_data[76][75] = 0;
        pixel_data[76][76] = 0;
        pixel_data[76][77] = 0;
        pixel_data[76][78] = 0;
        pixel_data[76][79] = 0;
        pixel_data[76][80] = 0;
        pixel_data[76][81] = 0;
        pixel_data[76][82] = 0;
        pixel_data[76][83] = 0;
        pixel_data[76][84] = 0;
        pixel_data[76][85] = 0;
        pixel_data[76][86] = 0;
        pixel_data[76][87] = 0;
        pixel_data[76][88] = 0;
        pixel_data[76][89] = 0;
        pixel_data[76][90] = 0;
        pixel_data[76][91] = 0;
        pixel_data[76][92] = 0;
        pixel_data[76][93] = 0;
        pixel_data[76][94] = 0;
        pixel_data[76][95] = 0;
        pixel_data[76][96] = 0;
        pixel_data[76][97] = 0;
        pixel_data[76][98] = 0;
        pixel_data[76][99] = 0; // y=76
        pixel_data[77][0] = 0;
        pixel_data[77][1] = 0;
        pixel_data[77][2] = 0;
        pixel_data[77][3] = 0;
        pixel_data[77][4] = 0;
        pixel_data[77][5] = 0;
        pixel_data[77][6] = 0;
        pixel_data[77][7] = 0;
        pixel_data[77][8] = 0;
        pixel_data[77][9] = 0;
        pixel_data[77][10] = 0;
        pixel_data[77][11] = 2;
        pixel_data[77][12] = 5;
        pixel_data[77][13] = 8;
        pixel_data[77][14] = 6;
        pixel_data[77][15] = 6;
        pixel_data[77][16] = 6;
        pixel_data[77][17] = 8;
        pixel_data[77][18] = 7;
        pixel_data[77][19] = 0;
        pixel_data[77][20] = 0;
        pixel_data[77][21] = 0;
        pixel_data[77][22] = 0;
        pixel_data[77][23] = 0;
        pixel_data[77][24] = 0;
        pixel_data[77][25] = 0;
        pixel_data[77][26] = 0;
        pixel_data[77][27] = 0;
        pixel_data[77][28] = 0;
        pixel_data[77][29] = 0;
        pixel_data[77][30] = 0;
        pixel_data[77][31] = 0;
        pixel_data[77][32] = 0;
        pixel_data[77][33] = 0;
        pixel_data[77][34] = 0;
        pixel_data[77][35] = 0;
        pixel_data[77][36] = 0;
        pixel_data[77][37] = 0;
        pixel_data[77][38] = 0;
        pixel_data[77][39] = 0;
        pixel_data[77][40] = 0;
        pixel_data[77][41] = 0;
        pixel_data[77][42] = 0;
        pixel_data[77][43] = 0;
        pixel_data[77][44] = 0;
        pixel_data[77][45] = 0;
        pixel_data[77][46] = 0;
        pixel_data[77][47] = 0;
        pixel_data[77][48] = 0;
        pixel_data[77][49] = 0;
        pixel_data[77][50] = 0;
        pixel_data[77][51] = 0;
        pixel_data[77][52] = 0;
        pixel_data[77][53] = 0;
        pixel_data[77][54] = 0;
        pixel_data[77][55] = 0;
        pixel_data[77][56] = 0;
        pixel_data[77][57] = 0;
        pixel_data[77][58] = 0;
        pixel_data[77][59] = 0;
        pixel_data[77][60] = 0;
        pixel_data[77][61] = 0;
        pixel_data[77][62] = 0;
        pixel_data[77][63] = 0;
        pixel_data[77][64] = 0;
        pixel_data[77][65] = 0;
        pixel_data[77][66] = 0;
        pixel_data[77][67] = 0;
        pixel_data[77][68] = 0;
        pixel_data[77][69] = 0;
        pixel_data[77][70] = 0;
        pixel_data[77][71] = 0;
        pixel_data[77][72] = 0;
        pixel_data[77][73] = 0;
        pixel_data[77][74] = 0;
        pixel_data[77][75] = 0;
        pixel_data[77][76] = 0;
        pixel_data[77][77] = 0;
        pixel_data[77][78] = 0;
        pixel_data[77][79] = 0;
        pixel_data[77][80] = 0;
        pixel_data[77][81] = 0;
        pixel_data[77][82] = 0;
        pixel_data[77][83] = 0;
        pixel_data[77][84] = 0;
        pixel_data[77][85] = 0;
        pixel_data[77][86] = 0;
        pixel_data[77][87] = 0;
        pixel_data[77][88] = 0;
        pixel_data[77][89] = 0;
        pixel_data[77][90] = 0;
        pixel_data[77][91] = 0;
        pixel_data[77][92] = 0;
        pixel_data[77][93] = 0;
        pixel_data[77][94] = 0;
        pixel_data[77][95] = 0;
        pixel_data[77][96] = 0;
        pixel_data[77][97] = 0;
        pixel_data[77][98] = 0;
        pixel_data[77][99] = 0; // y=77
        pixel_data[78][0] = 0;
        pixel_data[78][1] = 0;
        pixel_data[78][2] = 0;
        pixel_data[78][3] = 0;
        pixel_data[78][4] = 0;
        pixel_data[78][5] = 0;
        pixel_data[78][6] = 0;
        pixel_data[78][7] = 0;
        pixel_data[78][8] = 0;
        pixel_data[78][9] = 0;
        pixel_data[78][10] = 0;
        pixel_data[78][11] = 0;
        pixel_data[78][12] = 0;
        pixel_data[78][13] = 0;
        pixel_data[78][14] = 15;
        pixel_data[78][15] = 5;
        pixel_data[78][16] = 7;
        pixel_data[78][17] = 0;
        pixel_data[78][18] = 0;
        pixel_data[78][19] = 0;
        pixel_data[78][20] = 0;
        pixel_data[78][21] = 0;
        pixel_data[78][22] = 0;
        pixel_data[78][23] = 0;
        pixel_data[78][24] = 0;
        pixel_data[78][25] = 0;
        pixel_data[78][26] = 0;
        pixel_data[78][27] = 0;
        pixel_data[78][28] = 0;
        pixel_data[78][29] = 0;
        pixel_data[78][30] = 0;
        pixel_data[78][31] = 0;
        pixel_data[78][32] = 0;
        pixel_data[78][33] = 0;
        pixel_data[78][34] = 0;
        pixel_data[78][35] = 0;
        pixel_data[78][36] = 0;
        pixel_data[78][37] = 0;
        pixel_data[78][38] = 0;
        pixel_data[78][39] = 0;
        pixel_data[78][40] = 0;
        pixel_data[78][41] = 0;
        pixel_data[78][42] = 0;
        pixel_data[78][43] = 0;
        pixel_data[78][44] = 0;
        pixel_data[78][45] = 0;
        pixel_data[78][46] = 0;
        pixel_data[78][47] = 0;
        pixel_data[78][48] = 0;
        pixel_data[78][49] = 0;
        pixel_data[78][50] = 0;
        pixel_data[78][51] = 0;
        pixel_data[78][52] = 0;
        pixel_data[78][53] = 0;
        pixel_data[78][54] = 0;
        pixel_data[78][55] = 0;
        pixel_data[78][56] = 0;
        pixel_data[78][57] = 0;
        pixel_data[78][58] = 0;
        pixel_data[78][59] = 0;
        pixel_data[78][60] = 0;
        pixel_data[78][61] = 0;
        pixel_data[78][62] = 0;
        pixel_data[78][63] = 0;
        pixel_data[78][64] = 0;
        pixel_data[78][65] = 0;
        pixel_data[78][66] = 0;
        pixel_data[78][67] = 0;
        pixel_data[78][68] = 0;
        pixel_data[78][69] = 0;
        pixel_data[78][70] = 0;
        pixel_data[78][71] = 0;
        pixel_data[78][72] = 0;
        pixel_data[78][73] = 0;
        pixel_data[78][74] = 0;
        pixel_data[78][75] = 0;
        pixel_data[78][76] = 0;
        pixel_data[78][77] = 0;
        pixel_data[78][78] = 0;
        pixel_data[78][79] = 0;
        pixel_data[78][80] = 0;
        pixel_data[78][81] = 0;
        pixel_data[78][82] = 0;
        pixel_data[78][83] = 0;
        pixel_data[78][84] = 0;
        pixel_data[78][85] = 0;
        pixel_data[78][86] = 0;
        pixel_data[78][87] = 0;
        pixel_data[78][88] = 0;
        pixel_data[78][89] = 0;
        pixel_data[78][90] = 0;
        pixel_data[78][91] = 0;
        pixel_data[78][92] = 0;
        pixel_data[78][93] = 0;
        pixel_data[78][94] = 0;
        pixel_data[78][95] = 0;
        pixel_data[78][96] = 0;
        pixel_data[78][97] = 0;
        pixel_data[78][98] = 0;
        pixel_data[78][99] = 0; // y=78
        pixel_data[79][0] = 0;
        pixel_data[79][1] = 0;
        pixel_data[79][2] = 0;
        pixel_data[79][3] = 0;
        pixel_data[79][4] = 0;
        pixel_data[79][5] = 0;
        pixel_data[79][6] = 0;
        pixel_data[79][7] = 0;
        pixel_data[79][8] = 0;
        pixel_data[79][9] = 0;
        pixel_data[79][10] = 0;
        pixel_data[79][11] = 0;
        pixel_data[79][12] = 0;
        pixel_data[79][13] = 0;
        pixel_data[79][14] = 0;
        pixel_data[79][15] = 0;
        pixel_data[79][16] = 0;
        pixel_data[79][17] = 0;
        pixel_data[79][18] = 0;
        pixel_data[79][19] = 0;
        pixel_data[79][20] = 0;
        pixel_data[79][21] = 0;
        pixel_data[79][22] = 0;
        pixel_data[79][23] = 0;
        pixel_data[79][24] = 0;
        pixel_data[79][25] = 0;
        pixel_data[79][26] = 0;
        pixel_data[79][27] = 0;
        pixel_data[79][28] = 0;
        pixel_data[79][29] = 0;
        pixel_data[79][30] = 0;
        pixel_data[79][31] = 0;
        pixel_data[79][32] = 0;
        pixel_data[79][33] = 0;
        pixel_data[79][34] = 0;
        pixel_data[79][35] = 0;
        pixel_data[79][36] = 0;
        pixel_data[79][37] = 0;
        pixel_data[79][38] = 0;
        pixel_data[79][39] = 0;
        pixel_data[79][40] = 0;
        pixel_data[79][41] = 0;
        pixel_data[79][42] = 0;
        pixel_data[79][43] = 0;
        pixel_data[79][44] = 0;
        pixel_data[79][45] = 0;
        pixel_data[79][46] = 0;
        pixel_data[79][47] = 0;
        pixel_data[79][48] = 0;
        pixel_data[79][49] = 0;
        pixel_data[79][50] = 0;
        pixel_data[79][51] = 0;
        pixel_data[79][52] = 0;
        pixel_data[79][53] = 0;
        pixel_data[79][54] = 0;
        pixel_data[79][55] = 0;
        pixel_data[79][56] = 0;
        pixel_data[79][57] = 0;
        pixel_data[79][58] = 0;
        pixel_data[79][59] = 0;
        pixel_data[79][60] = 0;
        pixel_data[79][61] = 0;
        pixel_data[79][62] = 0;
        pixel_data[79][63] = 0;
        pixel_data[79][64] = 0;
        pixel_data[79][65] = 0;
        pixel_data[79][66] = 0;
        pixel_data[79][67] = 0;
        pixel_data[79][68] = 0;
        pixel_data[79][69] = 0;
        pixel_data[79][70] = 0;
        pixel_data[79][71] = 0;
        pixel_data[79][72] = 0;
        pixel_data[79][73] = 0;
        pixel_data[79][74] = 0;
        pixel_data[79][75] = 0;
        pixel_data[79][76] = 0;
        pixel_data[79][77] = 0;
        pixel_data[79][78] = 0;
        pixel_data[79][79] = 0;
        pixel_data[79][80] = 0;
        pixel_data[79][81] = 0;
        pixel_data[79][82] = 0;
        pixel_data[79][83] = 0;
        pixel_data[79][84] = 0;
        pixel_data[79][85] = 0;
        pixel_data[79][86] = 0;
        pixel_data[79][87] = 0;
        pixel_data[79][88] = 0;
        pixel_data[79][89] = 0;
        pixel_data[79][90] = 0;
        pixel_data[79][91] = 0;
        pixel_data[79][92] = 0;
        pixel_data[79][93] = 0;
        pixel_data[79][94] = 0;
        pixel_data[79][95] = 0;
        pixel_data[79][96] = 0;
        pixel_data[79][97] = 0;
        pixel_data[79][98] = 0;
        pixel_data[79][99] = 0; // y=79
        pixel_data[80][0] = 0;
        pixel_data[80][1] = 0;
        pixel_data[80][2] = 0;
        pixel_data[80][3] = 0;
        pixel_data[80][4] = 0;
        pixel_data[80][5] = 0;
        pixel_data[80][6] = 0;
        pixel_data[80][7] = 0;
        pixel_data[80][8] = 0;
        pixel_data[80][9] = 0;
        pixel_data[80][10] = 0;
        pixel_data[80][11] = 0;
        pixel_data[80][12] = 0;
        pixel_data[80][13] = 0;
        pixel_data[80][14] = 0;
        pixel_data[80][15] = 0;
        pixel_data[80][16] = 0;
        pixel_data[80][17] = 0;
        pixel_data[80][18] = 0;
        pixel_data[80][19] = 0;
        pixel_data[80][20] = 0;
        pixel_data[80][21] = 0;
        pixel_data[80][22] = 0;
        pixel_data[80][23] = 0;
        pixel_data[80][24] = 0;
        pixel_data[80][25] = 0;
        pixel_data[80][26] = 0;
        pixel_data[80][27] = 0;
        pixel_data[80][28] = 0;
        pixel_data[80][29] = 0;
        pixel_data[80][30] = 0;
        pixel_data[80][31] = 0;
        pixel_data[80][32] = 0;
        pixel_data[80][33] = 0;
        pixel_data[80][34] = 0;
        pixel_data[80][35] = 0;
        pixel_data[80][36] = 0;
        pixel_data[80][37] = 0;
        pixel_data[80][38] = 0;
        pixel_data[80][39] = 0;
        pixel_data[80][40] = 0;
        pixel_data[80][41] = 0;
        pixel_data[80][42] = 0;
        pixel_data[80][43] = 0;
        pixel_data[80][44] = 0;
        pixel_data[80][45] = 0;
        pixel_data[80][46] = 0;
        pixel_data[80][47] = 0;
        pixel_data[80][48] = 0;
        pixel_data[80][49] = 0;
        pixel_data[80][50] = 0;
        pixel_data[80][51] = 0;
        pixel_data[80][52] = 0;
        pixel_data[80][53] = 0;
        pixel_data[80][54] = 0;
        pixel_data[80][55] = 0;
        pixel_data[80][56] = 0;
        pixel_data[80][57] = 0;
        pixel_data[80][58] = 0;
        pixel_data[80][59] = 0;
        pixel_data[80][60] = 0;
        pixel_data[80][61] = 0;
        pixel_data[80][62] = 0;
        pixel_data[80][63] = 0;
        pixel_data[80][64] = 0;
        pixel_data[80][65] = 0;
        pixel_data[80][66] = 0;
        pixel_data[80][67] = 0;
        pixel_data[80][68] = 0;
        pixel_data[80][69] = 0;
        pixel_data[80][70] = 0;
        pixel_data[80][71] = 0;
        pixel_data[80][72] = 0;
        pixel_data[80][73] = 0;
        pixel_data[80][74] = 0;
        pixel_data[80][75] = 0;
        pixel_data[80][76] = 0;
        pixel_data[80][77] = 0;
        pixel_data[80][78] = 0;
        pixel_data[80][79] = 0;
        pixel_data[80][80] = 0;
        pixel_data[80][81] = 0;
        pixel_data[80][82] = 0;
        pixel_data[80][83] = 0;
        pixel_data[80][84] = 0;
        pixel_data[80][85] = 0;
        pixel_data[80][86] = 0;
        pixel_data[80][87] = 0;
        pixel_data[80][88] = 0;
        pixel_data[80][89] = 0;
        pixel_data[80][90] = 0;
        pixel_data[80][91] = 0;
        pixel_data[80][92] = 0;
        pixel_data[80][93] = 0;
        pixel_data[80][94] = 0;
        pixel_data[80][95] = 0;
        pixel_data[80][96] = 0;
        pixel_data[80][97] = 0;
        pixel_data[80][98] = 0;
        pixel_data[80][99] = 0; // y=80
        pixel_data[81][0] = 0;
        pixel_data[81][1] = 0;
        pixel_data[81][2] = 0;
        pixel_data[81][3] = 0;
        pixel_data[81][4] = 0;
        pixel_data[81][5] = 0;
        pixel_data[81][6] = 0;
        pixel_data[81][7] = 0;
        pixel_data[81][8] = 0;
        pixel_data[81][9] = 0;
        pixel_data[81][10] = 0;
        pixel_data[81][11] = 0;
        pixel_data[81][12] = 0;
        pixel_data[81][13] = 0;
        pixel_data[81][14] = 0;
        pixel_data[81][15] = 0;
        pixel_data[81][16] = 0;
        pixel_data[81][17] = 0;
        pixel_data[81][18] = 0;
        pixel_data[81][19] = 0;
        pixel_data[81][20] = 0;
        pixel_data[81][21] = 0;
        pixel_data[81][22] = 0;
        pixel_data[81][23] = 0;
        pixel_data[81][24] = 0;
        pixel_data[81][25] = 0;
        pixel_data[81][26] = 0;
        pixel_data[81][27] = 0;
        pixel_data[81][28] = 0;
        pixel_data[81][29] = 0;
        pixel_data[81][30] = 0;
        pixel_data[81][31] = 0;
        pixel_data[81][32] = 0;
        pixel_data[81][33] = 0;
        pixel_data[81][34] = 0;
        pixel_data[81][35] = 0;
        pixel_data[81][36] = 0;
        pixel_data[81][37] = 0;
        pixel_data[81][38] = 0;
        pixel_data[81][39] = 0;
        pixel_data[81][40] = 0;
        pixel_data[81][41] = 0;
        pixel_data[81][42] = 0;
        pixel_data[81][43] = 0;
        pixel_data[81][44] = 0;
        pixel_data[81][45] = 0;
        pixel_data[81][46] = 0;
        pixel_data[81][47] = 0;
        pixel_data[81][48] = 0;
        pixel_data[81][49] = 0;
        pixel_data[81][50] = 0;
        pixel_data[81][51] = 0;
        pixel_data[81][52] = 0;
        pixel_data[81][53] = 0;
        pixel_data[81][54] = 0;
        pixel_data[81][55] = 0;
        pixel_data[81][56] = 0;
        pixel_data[81][57] = 0;
        pixel_data[81][58] = 0;
        pixel_data[81][59] = 0;
        pixel_data[81][60] = 0;
        pixel_data[81][61] = 0;
        pixel_data[81][62] = 0;
        pixel_data[81][63] = 0;
        pixel_data[81][64] = 0;
        pixel_data[81][65] = 0;
        pixel_data[81][66] = 0;
        pixel_data[81][67] = 0;
        pixel_data[81][68] = 0;
        pixel_data[81][69] = 0;
        pixel_data[81][70] = 0;
        pixel_data[81][71] = 0;
        pixel_data[81][72] = 0;
        pixel_data[81][73] = 0;
        pixel_data[81][74] = 0;
        pixel_data[81][75] = 0;
        pixel_data[81][76] = 0;
        pixel_data[81][77] = 0;
        pixel_data[81][78] = 0;
        pixel_data[81][79] = 0;
        pixel_data[81][80] = 0;
        pixel_data[81][81] = 0;
        pixel_data[81][82] = 0;
        pixel_data[81][83] = 0;
        pixel_data[81][84] = 0;
        pixel_data[81][85] = 0;
        pixel_data[81][86] = 0;
        pixel_data[81][87] = 0;
        pixel_data[81][88] = 0;
        pixel_data[81][89] = 0;
        pixel_data[81][90] = 0;
        pixel_data[81][91] = 0;
        pixel_data[81][92] = 0;
        pixel_data[81][93] = 0;
        pixel_data[81][94] = 0;
        pixel_data[81][95] = 0;
        pixel_data[81][96] = 0;
        pixel_data[81][97] = 0;
        pixel_data[81][98] = 0;
        pixel_data[81][99] = 0; // y=81
        pixel_data[82][0] = 0;
        pixel_data[82][1] = 0;
        pixel_data[82][2] = 0;
        pixel_data[82][3] = 0;
        pixel_data[82][4] = 0;
        pixel_data[82][5] = 0;
        pixel_data[82][6] = 0;
        pixel_data[82][7] = 0;
        pixel_data[82][8] = 0;
        pixel_data[82][9] = 0;
        pixel_data[82][10] = 0;
        pixel_data[82][11] = 0;
        pixel_data[82][12] = 0;
        pixel_data[82][13] = 0;
        pixel_data[82][14] = 0;
        pixel_data[82][15] = 0;
        pixel_data[82][16] = 0;
        pixel_data[82][17] = 0;
        pixel_data[82][18] = 0;
        pixel_data[82][19] = 0;
        pixel_data[82][20] = 0;
        pixel_data[82][21] = 0;
        pixel_data[82][22] = 0;
        pixel_data[82][23] = 0;
        pixel_data[82][24] = 0;
        pixel_data[82][25] = 0;
        pixel_data[82][26] = 0;
        pixel_data[82][27] = 0;
        pixel_data[82][28] = 0;
        pixel_data[82][29] = 0;
        pixel_data[82][30] = 0;
        pixel_data[82][31] = 0;
        pixel_data[82][32] = 0;
        pixel_data[82][33] = 0;
        pixel_data[82][34] = 0;
        pixel_data[82][35] = 0;
        pixel_data[82][36] = 0;
        pixel_data[82][37] = 0;
        pixel_data[82][38] = 0;
        pixel_data[82][39] = 0;
        pixel_data[82][40] = 0;
        pixel_data[82][41] = 0;
        pixel_data[82][42] = 0;
        pixel_data[82][43] = 0;
        pixel_data[82][44] = 0;
        pixel_data[82][45] = 0;
        pixel_data[82][46] = 0;
        pixel_data[82][47] = 0;
        pixel_data[82][48] = 0;
        pixel_data[82][49] = 0;
        pixel_data[82][50] = 0;
        pixel_data[82][51] = 0;
        pixel_data[82][52] = 0;
        pixel_data[82][53] = 0;
        pixel_data[82][54] = 0;
        pixel_data[82][55] = 0;
        pixel_data[82][56] = 0;
        pixel_data[82][57] = 0;
        pixel_data[82][58] = 0;
        pixel_data[82][59] = 0;
        pixel_data[82][60] = 0;
        pixel_data[82][61] = 0;
        pixel_data[82][62] = 0;
        pixel_data[82][63] = 0;
        pixel_data[82][64] = 0;
        pixel_data[82][65] = 0;
        pixel_data[82][66] = 0;
        pixel_data[82][67] = 0;
        pixel_data[82][68] = 0;
        pixel_data[82][69] = 0;
        pixel_data[82][70] = 0;
        pixel_data[82][71] = 0;
        pixel_data[82][72] = 0;
        pixel_data[82][73] = 0;
        pixel_data[82][74] = 0;
        pixel_data[82][75] = 0;
        pixel_data[82][76] = 0;
        pixel_data[82][77] = 0;
        pixel_data[82][78] = 0;
        pixel_data[82][79] = 0;
        pixel_data[82][80] = 0;
        pixel_data[82][81] = 0;
        pixel_data[82][82] = 0;
        pixel_data[82][83] = 0;
        pixel_data[82][84] = 0;
        pixel_data[82][85] = 0;
        pixel_data[82][86] = 0;
        pixel_data[82][87] = 0;
        pixel_data[82][88] = 0;
        pixel_data[82][89] = 0;
        pixel_data[82][90] = 0;
        pixel_data[82][91] = 0;
        pixel_data[82][92] = 0;
        pixel_data[82][93] = 0;
        pixel_data[82][94] = 0;
        pixel_data[82][95] = 0;
        pixel_data[82][96] = 0;
        pixel_data[82][97] = 0;
        pixel_data[82][98] = 0;
        pixel_data[82][99] = 0; // y=82
        pixel_data[83][0] = 0;
        pixel_data[83][1] = 0;
        pixel_data[83][2] = 0;
        pixel_data[83][3] = 0;
        pixel_data[83][4] = 0;
        pixel_data[83][5] = 0;
        pixel_data[83][6] = 0;
        pixel_data[83][7] = 0;
        pixel_data[83][8] = 0;
        pixel_data[83][9] = 0;
        pixel_data[83][10] = 0;
        pixel_data[83][11] = 0;
        pixel_data[83][12] = 0;
        pixel_data[83][13] = 0;
        pixel_data[83][14] = 0;
        pixel_data[83][15] = 0;
        pixel_data[83][16] = 0;
        pixel_data[83][17] = 0;
        pixel_data[83][18] = 0;
        pixel_data[83][19] = 0;
        pixel_data[83][20] = 0;
        pixel_data[83][21] = 0;
        pixel_data[83][22] = 0;
        pixel_data[83][23] = 0;
        pixel_data[83][24] = 0;
        pixel_data[83][25] = 0;
        pixel_data[83][26] = 0;
        pixel_data[83][27] = 0;
        pixel_data[83][28] = 0;
        pixel_data[83][29] = 0;
        pixel_data[83][30] = 0;
        pixel_data[83][31] = 0;
        pixel_data[83][32] = 0;
        pixel_data[83][33] = 0;
        pixel_data[83][34] = 0;
        pixel_data[83][35] = 0;
        pixel_data[83][36] = 0;
        pixel_data[83][37] = 0;
        pixel_data[83][38] = 0;
        pixel_data[83][39] = 0;
        pixel_data[83][40] = 0;
        pixel_data[83][41] = 0;
        pixel_data[83][42] = 0;
        pixel_data[83][43] = 0;
        pixel_data[83][44] = 0;
        pixel_data[83][45] = 0;
        pixel_data[83][46] = 0;
        pixel_data[83][47] = 0;
        pixel_data[83][48] = 0;
        pixel_data[83][49] = 0;
        pixel_data[83][50] = 0;
        pixel_data[83][51] = 0;
        pixel_data[83][52] = 0;
        pixel_data[83][53] = 0;
        pixel_data[83][54] = 0;
        pixel_data[83][55] = 0;
        pixel_data[83][56] = 0;
        pixel_data[83][57] = 0;
        pixel_data[83][58] = 0;
        pixel_data[83][59] = 0;
        pixel_data[83][60] = 0;
        pixel_data[83][61] = 0;
        pixel_data[83][62] = 0;
        pixel_data[83][63] = 0;
        pixel_data[83][64] = 0;
        pixel_data[83][65] = 0;
        pixel_data[83][66] = 0;
        pixel_data[83][67] = 0;
        pixel_data[83][68] = 0;
        pixel_data[83][69] = 0;
        pixel_data[83][70] = 0;
        pixel_data[83][71] = 0;
        pixel_data[83][72] = 0;
        pixel_data[83][73] = 0;
        pixel_data[83][74] = 0;
        pixel_data[83][75] = 0;
        pixel_data[83][76] = 0;
        pixel_data[83][77] = 0;
        pixel_data[83][78] = 0;
        pixel_data[83][79] = 0;
        pixel_data[83][80] = 0;
        pixel_data[83][81] = 0;
        pixel_data[83][82] = 0;
        pixel_data[83][83] = 0;
        pixel_data[83][84] = 0;
        pixel_data[83][85] = 0;
        pixel_data[83][86] = 0;
        pixel_data[83][87] = 0;
        pixel_data[83][88] = 0;
        pixel_data[83][89] = 0;
        pixel_data[83][90] = 0;
        pixel_data[83][91] = 0;
        pixel_data[83][92] = 0;
        pixel_data[83][93] = 0;
        pixel_data[83][94] = 0;
        pixel_data[83][95] = 0;
        pixel_data[83][96] = 0;
        pixel_data[83][97] = 0;
        pixel_data[83][98] = 0;
        pixel_data[83][99] = 0; // y=83
        pixel_data[84][0] = 0;
        pixel_data[84][1] = 0;
        pixel_data[84][2] = 0;
        pixel_data[84][3] = 0;
        pixel_data[84][4] = 0;
        pixel_data[84][5] = 0;
        pixel_data[84][6] = 0;
        pixel_data[84][7] = 0;
        pixel_data[84][8] = 0;
        pixel_data[84][9] = 0;
        pixel_data[84][10] = 0;
        pixel_data[84][11] = 0;
        pixel_data[84][12] = 0;
        pixel_data[84][13] = 0;
        pixel_data[84][14] = 0;
        pixel_data[84][15] = 0;
        pixel_data[84][16] = 0;
        pixel_data[84][17] = 0;
        pixel_data[84][18] = 0;
        pixel_data[84][19] = 0;
        pixel_data[84][20] = 0;
        pixel_data[84][21] = 0;
        pixel_data[84][22] = 0;
        pixel_data[84][23] = 0;
        pixel_data[84][24] = 0;
        pixel_data[84][25] = 0;
        pixel_data[84][26] = 0;
        pixel_data[84][27] = 0;
        pixel_data[84][28] = 0;
        pixel_data[84][29] = 0;
        pixel_data[84][30] = 0;
        pixel_data[84][31] = 0;
        pixel_data[84][32] = 0;
        pixel_data[84][33] = 0;
        pixel_data[84][34] = 0;
        pixel_data[84][35] = 0;
        pixel_data[84][36] = 0;
        pixel_data[84][37] = 0;
        pixel_data[84][38] = 0;
        pixel_data[84][39] = 0;
        pixel_data[84][40] = 0;
        pixel_data[84][41] = 0;
        pixel_data[84][42] = 0;
        pixel_data[84][43] = 0;
        pixel_data[84][44] = 0;
        pixel_data[84][45] = 0;
        pixel_data[84][46] = 0;
        pixel_data[84][47] = 0;
        pixel_data[84][48] = 0;
        pixel_data[84][49] = 0;
        pixel_data[84][50] = 0;
        pixel_data[84][51] = 0;
        pixel_data[84][52] = 0;
        pixel_data[84][53] = 0;
        pixel_data[84][54] = 0;
        pixel_data[84][55] = 0;
        pixel_data[84][56] = 0;
        pixel_data[84][57] = 0;
        pixel_data[84][58] = 0;
        pixel_data[84][59] = 0;
        pixel_data[84][60] = 0;
        pixel_data[84][61] = 0;
        pixel_data[84][62] = 0;
        pixel_data[84][63] = 0;
        pixel_data[84][64] = 0;
        pixel_data[84][65] = 0;
        pixel_data[84][66] = 0;
        pixel_data[84][67] = 0;
        pixel_data[84][68] = 0;
        pixel_data[84][69] = 0;
        pixel_data[84][70] = 0;
        pixel_data[84][71] = 0;
        pixel_data[84][72] = 0;
        pixel_data[84][73] = 0;
        pixel_data[84][74] = 0;
        pixel_data[84][75] = 0;
        pixel_data[84][76] = 0;
        pixel_data[84][77] = 0;
        pixel_data[84][78] = 0;
        pixel_data[84][79] = 0;
        pixel_data[84][80] = 0;
        pixel_data[84][81] = 0;
        pixel_data[84][82] = 0;
        pixel_data[84][83] = 0;
        pixel_data[84][84] = 0;
        pixel_data[84][85] = 0;
        pixel_data[84][86] = 0;
        pixel_data[84][87] = 0;
        pixel_data[84][88] = 0;
        pixel_data[84][89] = 0;
        pixel_data[84][90] = 0;
        pixel_data[84][91] = 0;
        pixel_data[84][92] = 0;
        pixel_data[84][93] = 0;
        pixel_data[84][94] = 0;
        pixel_data[84][95] = 0;
        pixel_data[84][96] = 0;
        pixel_data[84][97] = 0;
        pixel_data[84][98] = 0;
        pixel_data[84][99] = 0; // y=84
        pixel_data[85][0] = 0;
        pixel_data[85][1] = 0;
        pixel_data[85][2] = 0;
        pixel_data[85][3] = 0;
        pixel_data[85][4] = 0;
        pixel_data[85][5] = 0;
        pixel_data[85][6] = 0;
        pixel_data[85][7] = 0;
        pixel_data[85][8] = 0;
        pixel_data[85][9] = 0;
        pixel_data[85][10] = 0;
        pixel_data[85][11] = 0;
        pixel_data[85][12] = 0;
        pixel_data[85][13] = 0;
        pixel_data[85][14] = 0;
        pixel_data[85][15] = 0;
        pixel_data[85][16] = 0;
        pixel_data[85][17] = 0;
        pixel_data[85][18] = 0;
        pixel_data[85][19] = 0;
        pixel_data[85][20] = 0;
        pixel_data[85][21] = 0;
        pixel_data[85][22] = 0;
        pixel_data[85][23] = 0;
        pixel_data[85][24] = 0;
        pixel_data[85][25] = 0;
        pixel_data[85][26] = 0;
        pixel_data[85][27] = 0;
        pixel_data[85][28] = 0;
        pixel_data[85][29] = 0;
        pixel_data[85][30] = 0;
        pixel_data[85][31] = 0;
        pixel_data[85][32] = 0;
        pixel_data[85][33] = 0;
        pixel_data[85][34] = 0;
        pixel_data[85][35] = 0;
        pixel_data[85][36] = 0;
        pixel_data[85][37] = 0;
        pixel_data[85][38] = 0;
        pixel_data[85][39] = 0;
        pixel_data[85][40] = 0;
        pixel_data[85][41] = 0;
        pixel_data[85][42] = 0;
        pixel_data[85][43] = 0;
        pixel_data[85][44] = 0;
        pixel_data[85][45] = 0;
        pixel_data[85][46] = 0;
        pixel_data[85][47] = 0;
        pixel_data[85][48] = 0;
        pixel_data[85][49] = 0;
        pixel_data[85][50] = 0;
        pixel_data[85][51] = 0;
        pixel_data[85][52] = 0;
        pixel_data[85][53] = 0;
        pixel_data[85][54] = 0;
        pixel_data[85][55] = 0;
        pixel_data[85][56] = 0;
        pixel_data[85][57] = 0;
        pixel_data[85][58] = 0;
        pixel_data[85][59] = 0;
        pixel_data[85][60] = 0;
        pixel_data[85][61] = 0;
        pixel_data[85][62] = 0;
        pixel_data[85][63] = 0;
        pixel_data[85][64] = 0;
        pixel_data[85][65] = 0;
        pixel_data[85][66] = 0;
        pixel_data[85][67] = 0;
        pixel_data[85][68] = 0;
        pixel_data[85][69] = 0;
        pixel_data[85][70] = 0;
        pixel_data[85][71] = 0;
        pixel_data[85][72] = 0;
        pixel_data[85][73] = 0;
        pixel_data[85][74] = 0;
        pixel_data[85][75] = 0;
        pixel_data[85][76] = 0;
        pixel_data[85][77] = 0;
        pixel_data[85][78] = 0;
        pixel_data[85][79] = 0;
        pixel_data[85][80] = 0;
        pixel_data[85][81] = 0;
        pixel_data[85][82] = 0;
        pixel_data[85][83] = 0;
        pixel_data[85][84] = 0;
        pixel_data[85][85] = 0;
        pixel_data[85][86] = 0;
        pixel_data[85][87] = 0;
        pixel_data[85][88] = 0;
        pixel_data[85][89] = 0;
        pixel_data[85][90] = 0;
        pixel_data[85][91] = 0;
        pixel_data[85][92] = 0;
        pixel_data[85][93] = 0;
        pixel_data[85][94] = 0;
        pixel_data[85][95] = 0;
        pixel_data[85][96] = 0;
        pixel_data[85][97] = 0;
        pixel_data[85][98] = 0;
        pixel_data[85][99] = 0; // y=85
        pixel_data[86][0] = 0;
        pixel_data[86][1] = 0;
        pixel_data[86][2] = 0;
        pixel_data[86][3] = 0;
        pixel_data[86][4] = 0;
        pixel_data[86][5] = 0;
        pixel_data[86][6] = 0;
        pixel_data[86][7] = 0;
        pixel_data[86][8] = 0;
        pixel_data[86][9] = 0;
        pixel_data[86][10] = 0;
        pixel_data[86][11] = 0;
        pixel_data[86][12] = 0;
        pixel_data[86][13] = 0;
        pixel_data[86][14] = 0;
        pixel_data[86][15] = 0;
        pixel_data[86][16] = 0;
        pixel_data[86][17] = 0;
        pixel_data[86][18] = 0;
        pixel_data[86][19] = 0;
        pixel_data[86][20] = 0;
        pixel_data[86][21] = 0;
        pixel_data[86][22] = 0;
        pixel_data[86][23] = 0;
        pixel_data[86][24] = 0;
        pixel_data[86][25] = 0;
        pixel_data[86][26] = 0;
        pixel_data[86][27] = 0;
        pixel_data[86][28] = 0;
        pixel_data[86][29] = 0;
        pixel_data[86][30] = 0;
        pixel_data[86][31] = 0;
        pixel_data[86][32] = 0;
        pixel_data[86][33] = 0;
        pixel_data[86][34] = 0;
        pixel_data[86][35] = 0;
        pixel_data[86][36] = 0;
        pixel_data[86][37] = 0;
        pixel_data[86][38] = 0;
        pixel_data[86][39] = 0;
        pixel_data[86][40] = 0;
        pixel_data[86][41] = 0;
        pixel_data[86][42] = 0;
        pixel_data[86][43] = 0;
        pixel_data[86][44] = 0;
        pixel_data[86][45] = 0;
        pixel_data[86][46] = 0;
        pixel_data[86][47] = 0;
        pixel_data[86][48] = 0;
        pixel_data[86][49] = 0;
        pixel_data[86][50] = 0;
        pixel_data[86][51] = 0;
        pixel_data[86][52] = 0;
        pixel_data[86][53] = 0;
        pixel_data[86][54] = 0;
        pixel_data[86][55] = 0;
        pixel_data[86][56] = 0;
        pixel_data[86][57] = 0;
        pixel_data[86][58] = 0;
        pixel_data[86][59] = 0;
        pixel_data[86][60] = 0;
        pixel_data[86][61] = 0;
        pixel_data[86][62] = 0;
        pixel_data[86][63] = 0;
        pixel_data[86][64] = 0;
        pixel_data[86][65] = 0;
        pixel_data[86][66] = 0;
        pixel_data[86][67] = 0;
        pixel_data[86][68] = 0;
        pixel_data[86][69] = 0;
        pixel_data[86][70] = 0;
        pixel_data[86][71] = 0;
        pixel_data[86][72] = 0;
        pixel_data[86][73] = 0;
        pixel_data[86][74] = 0;
        pixel_data[86][75] = 0;
        pixel_data[86][76] = 0;
        pixel_data[86][77] = 0;
        pixel_data[86][78] = 0;
        pixel_data[86][79] = 0;
        pixel_data[86][80] = 0;
        pixel_data[86][81] = 0;
        pixel_data[86][82] = 0;
        pixel_data[86][83] = 0;
        pixel_data[86][84] = 0;
        pixel_data[86][85] = 0;
        pixel_data[86][86] = 0;
        pixel_data[86][87] = 0;
        pixel_data[86][88] = 0;
        pixel_data[86][89] = 0;
        pixel_data[86][90] = 0;
        pixel_data[86][91] = 0;
        pixel_data[86][92] = 0;
        pixel_data[86][93] = 0;
        pixel_data[86][94] = 0;
        pixel_data[86][95] = 0;
        pixel_data[86][96] = 0;
        pixel_data[86][97] = 0;
        pixel_data[86][98] = 0;
        pixel_data[86][99] = 0; // y=86
        pixel_data[87][0] = 0;
        pixel_data[87][1] = 0;
        pixel_data[87][2] = 0;
        pixel_data[87][3] = 0;
        pixel_data[87][4] = 0;
        pixel_data[87][5] = 0;
        pixel_data[87][6] = 0;
        pixel_data[87][7] = 0;
        pixel_data[87][8] = 0;
        pixel_data[87][9] = 0;
        pixel_data[87][10] = 0;
        pixel_data[87][11] = 0;
        pixel_data[87][12] = 0;
        pixel_data[87][13] = 0;
        pixel_data[87][14] = 0;
        pixel_data[87][15] = 0;
        pixel_data[87][16] = 0;
        pixel_data[87][17] = 0;
        pixel_data[87][18] = 0;
        pixel_data[87][19] = 0;
        pixel_data[87][20] = 0;
        pixel_data[87][21] = 0;
        pixel_data[87][22] = 0;
        pixel_data[87][23] = 0;
        pixel_data[87][24] = 0;
        pixel_data[87][25] = 0;
        pixel_data[87][26] = 0;
        pixel_data[87][27] = 0;
        pixel_data[87][28] = 0;
        pixel_data[87][29] = 0;
        pixel_data[87][30] = 0;
        pixel_data[87][31] = 0;
        pixel_data[87][32] = 0;
        pixel_data[87][33] = 0;
        pixel_data[87][34] = 0;
        pixel_data[87][35] = 0;
        pixel_data[87][36] = 0;
        pixel_data[87][37] = 0;
        pixel_data[87][38] = 0;
        pixel_data[87][39] = 0;
        pixel_data[87][40] = 0;
        pixel_data[87][41] = 0;
        pixel_data[87][42] = 0;
        pixel_data[87][43] = 0;
        pixel_data[87][44] = 0;
        pixel_data[87][45] = 0;
        pixel_data[87][46] = 0;
        pixel_data[87][47] = 0;
        pixel_data[87][48] = 0;
        pixel_data[87][49] = 0;
        pixel_data[87][50] = 0;
        pixel_data[87][51] = 0;
        pixel_data[87][52] = 0;
        pixel_data[87][53] = 0;
        pixel_data[87][54] = 0;
        pixel_data[87][55] = 0;
        pixel_data[87][56] = 0;
        pixel_data[87][57] = 0;
        pixel_data[87][58] = 0;
        pixel_data[87][59] = 0;
        pixel_data[87][60] = 0;
        pixel_data[87][61] = 0;
        pixel_data[87][62] = 0;
        pixel_data[87][63] = 0;
        pixel_data[87][64] = 0;
        pixel_data[87][65] = 0;
        pixel_data[87][66] = 0;
        pixel_data[87][67] = 0;
        pixel_data[87][68] = 0;
        pixel_data[87][69] = 0;
        pixel_data[87][70] = 0;
        pixel_data[87][71] = 0;
        pixel_data[87][72] = 0;
        pixel_data[87][73] = 0;
        pixel_data[87][74] = 0;
        pixel_data[87][75] = 0;
        pixel_data[87][76] = 0;
        pixel_data[87][77] = 0;
        pixel_data[87][78] = 0;
        pixel_data[87][79] = 0;
        pixel_data[87][80] = 0;
        pixel_data[87][81] = 0;
        pixel_data[87][82] = 0;
        pixel_data[87][83] = 0;
        pixel_data[87][84] = 0;
        pixel_data[87][85] = 0;
        pixel_data[87][86] = 0;
        pixel_data[87][87] = 0;
        pixel_data[87][88] = 0;
        pixel_data[87][89] = 0;
        pixel_data[87][90] = 0;
        pixel_data[87][91] = 0;
        pixel_data[87][92] = 0;
        pixel_data[87][93] = 0;
        pixel_data[87][94] = 0;
        pixel_data[87][95] = 0;
        pixel_data[87][96] = 0;
        pixel_data[87][97] = 0;
        pixel_data[87][98] = 0;
        pixel_data[87][99] = 0; // y=87
        pixel_data[88][0] = 0;
        pixel_data[88][1] = 0;
        pixel_data[88][2] = 0;
        pixel_data[88][3] = 0;
        pixel_data[88][4] = 0;
        pixel_data[88][5] = 0;
        pixel_data[88][6] = 0;
        pixel_data[88][7] = 0;
        pixel_data[88][8] = 0;
        pixel_data[88][9] = 0;
        pixel_data[88][10] = 0;
        pixel_data[88][11] = 0;
        pixel_data[88][12] = 0;
        pixel_data[88][13] = 0;
        pixel_data[88][14] = 0;
        pixel_data[88][15] = 0;
        pixel_data[88][16] = 0;
        pixel_data[88][17] = 0;
        pixel_data[88][18] = 0;
        pixel_data[88][19] = 0;
        pixel_data[88][20] = 0;
        pixel_data[88][21] = 0;
        pixel_data[88][22] = 0;
        pixel_data[88][23] = 0;
        pixel_data[88][24] = 0;
        pixel_data[88][25] = 0;
        pixel_data[88][26] = 0;
        pixel_data[88][27] = 0;
        pixel_data[88][28] = 0;
        pixel_data[88][29] = 0;
        pixel_data[88][30] = 0;
        pixel_data[88][31] = 0;
        pixel_data[88][32] = 0;
        pixel_data[88][33] = 0;
        pixel_data[88][34] = 0;
        pixel_data[88][35] = 0;
        pixel_data[88][36] = 0;
        pixel_data[88][37] = 0;
        pixel_data[88][38] = 0;
        pixel_data[88][39] = 0;
        pixel_data[88][40] = 0;
        pixel_data[88][41] = 0;
        pixel_data[88][42] = 0;
        pixel_data[88][43] = 0;
        pixel_data[88][44] = 0;
        pixel_data[88][45] = 0;
        pixel_data[88][46] = 0;
        pixel_data[88][47] = 0;
        pixel_data[88][48] = 0;
        pixel_data[88][49] = 0;
        pixel_data[88][50] = 0;
        pixel_data[88][51] = 0;
        pixel_data[88][52] = 0;
        pixel_data[88][53] = 0;
        pixel_data[88][54] = 0;
        pixel_data[88][55] = 0;
        pixel_data[88][56] = 0;
        pixel_data[88][57] = 0;
        pixel_data[88][58] = 0;
        pixel_data[88][59] = 0;
        pixel_data[88][60] = 0;
        pixel_data[88][61] = 0;
        pixel_data[88][62] = 0;
        pixel_data[88][63] = 0;
        pixel_data[88][64] = 0;
        pixel_data[88][65] = 0;
        pixel_data[88][66] = 0;
        pixel_data[88][67] = 0;
        pixel_data[88][68] = 0;
        pixel_data[88][69] = 0;
        pixel_data[88][70] = 0;
        pixel_data[88][71] = 0;
        pixel_data[88][72] = 0;
        pixel_data[88][73] = 0;
        pixel_data[88][74] = 0;
        pixel_data[88][75] = 0;
        pixel_data[88][76] = 0;
        pixel_data[88][77] = 0;
        pixel_data[88][78] = 0;
        pixel_data[88][79] = 0;
        pixel_data[88][80] = 0;
        pixel_data[88][81] = 0;
        pixel_data[88][82] = 0;
        pixel_data[88][83] = 0;
        pixel_data[88][84] = 0;
        pixel_data[88][85] = 0;
        pixel_data[88][86] = 0;
        pixel_data[88][87] = 0;
        pixel_data[88][88] = 0;
        pixel_data[88][89] = 0;
        pixel_data[88][90] = 0;
        pixel_data[88][91] = 0;
        pixel_data[88][92] = 0;
        pixel_data[88][93] = 0;
        pixel_data[88][94] = 0;
        pixel_data[88][95] = 0;
        pixel_data[88][96] = 0;
        pixel_data[88][97] = 0;
        pixel_data[88][98] = 0;
        pixel_data[88][99] = 0; // y=88
        pixel_data[89][0] = 0;
        pixel_data[89][1] = 0;
        pixel_data[89][2] = 0;
        pixel_data[89][3] = 0;
        pixel_data[89][4] = 0;
        pixel_data[89][5] = 0;
        pixel_data[89][6] = 0;
        pixel_data[89][7] = 0;
        pixel_data[89][8] = 0;
        pixel_data[89][9] = 0;
        pixel_data[89][10] = 0;
        pixel_data[89][11] = 0;
        pixel_data[89][12] = 0;
        pixel_data[89][13] = 0;
        pixel_data[89][14] = 0;
        pixel_data[89][15] = 0;
        pixel_data[89][16] = 0;
        pixel_data[89][17] = 0;
        pixel_data[89][18] = 0;
        pixel_data[89][19] = 0;
        pixel_data[89][20] = 0;
        pixel_data[89][21] = 0;
        pixel_data[89][22] = 0;
        pixel_data[89][23] = 0;
        pixel_data[89][24] = 0;
        pixel_data[89][25] = 0;
        pixel_data[89][26] = 0;
        pixel_data[89][27] = 0;
        pixel_data[89][28] = 0;
        pixel_data[89][29] = 0;
        pixel_data[89][30] = 0;
        pixel_data[89][31] = 0;
        pixel_data[89][32] = 0;
        pixel_data[89][33] = 0;
        pixel_data[89][34] = 0;
        pixel_data[89][35] = 0;
        pixel_data[89][36] = 0;
        pixel_data[89][37] = 0;
        pixel_data[89][38] = 0;
        pixel_data[89][39] = 0;
        pixel_data[89][40] = 0;
        pixel_data[89][41] = 0;
        pixel_data[89][42] = 0;
        pixel_data[89][43] = 0;
        pixel_data[89][44] = 0;
        pixel_data[89][45] = 0;
        pixel_data[89][46] = 0;
        pixel_data[89][47] = 0;
        pixel_data[89][48] = 0;
        pixel_data[89][49] = 0;
        pixel_data[89][50] = 0;
        pixel_data[89][51] = 0;
        pixel_data[89][52] = 0;
        pixel_data[89][53] = 0;
        pixel_data[89][54] = 0;
        pixel_data[89][55] = 0;
        pixel_data[89][56] = 0;
        pixel_data[89][57] = 0;
        pixel_data[89][58] = 0;
        pixel_data[89][59] = 0;
        pixel_data[89][60] = 0;
        pixel_data[89][61] = 0;
        pixel_data[89][62] = 0;
        pixel_data[89][63] = 0;
        pixel_data[89][64] = 0;
        pixel_data[89][65] = 0;
        pixel_data[89][66] = 0;
        pixel_data[89][67] = 0;
        pixel_data[89][68] = 0;
        pixel_data[89][69] = 0;
        pixel_data[89][70] = 0;
        pixel_data[89][71] = 0;
        pixel_data[89][72] = 0;
        pixel_data[89][73] = 0;
        pixel_data[89][74] = 0;
        pixel_data[89][75] = 0;
        pixel_data[89][76] = 0;
        pixel_data[89][77] = 0;
        pixel_data[89][78] = 0;
        pixel_data[89][79] = 0;
        pixel_data[89][80] = 0;
        pixel_data[89][81] = 0;
        pixel_data[89][82] = 0;
        pixel_data[89][83] = 0;
        pixel_data[89][84] = 0;
        pixel_data[89][85] = 0;
        pixel_data[89][86] = 0;
        pixel_data[89][87] = 0;
        pixel_data[89][88] = 0;
        pixel_data[89][89] = 0;
        pixel_data[89][90] = 0;
        pixel_data[89][91] = 0;
        pixel_data[89][92] = 0;
        pixel_data[89][93] = 0;
        pixel_data[89][94] = 0;
        pixel_data[89][95] = 0;
        pixel_data[89][96] = 0;
        pixel_data[89][97] = 0;
        pixel_data[89][98] = 0;
        pixel_data[89][99] = 0; // y=89
        pixel_data[90][0] = 0;
        pixel_data[90][1] = 0;
        pixel_data[90][2] = 0;
        pixel_data[90][3] = 0;
        pixel_data[90][4] = 0;
        pixel_data[90][5] = 0;
        pixel_data[90][6] = 0;
        pixel_data[90][7] = 0;
        pixel_data[90][8] = 0;
        pixel_data[90][9] = 0;
        pixel_data[90][10] = 0;
        pixel_data[90][11] = 0;
        pixel_data[90][12] = 0;
        pixel_data[90][13] = 0;
        pixel_data[90][14] = 0;
        pixel_data[90][15] = 0;
        pixel_data[90][16] = 0;
        pixel_data[90][17] = 0;
        pixel_data[90][18] = 0;
        pixel_data[90][19] = 0;
        pixel_data[90][20] = 0;
        pixel_data[90][21] = 0;
        pixel_data[90][22] = 0;
        pixel_data[90][23] = 0;
        pixel_data[90][24] = 0;
        pixel_data[90][25] = 0;
        pixel_data[90][26] = 0;
        pixel_data[90][27] = 0;
        pixel_data[90][28] = 0;
        pixel_data[90][29] = 0;
        pixel_data[90][30] = 0;
        pixel_data[90][31] = 0;
        pixel_data[90][32] = 0;
        pixel_data[90][33] = 0;
        pixel_data[90][34] = 0;
        pixel_data[90][35] = 0;
        pixel_data[90][36] = 0;
        pixel_data[90][37] = 0;
        pixel_data[90][38] = 0;
        pixel_data[90][39] = 0;
        pixel_data[90][40] = 0;
        pixel_data[90][41] = 0;
        pixel_data[90][42] = 0;
        pixel_data[90][43] = 0;
        pixel_data[90][44] = 0;
        pixel_data[90][45] = 0;
        pixel_data[90][46] = 0;
        pixel_data[90][47] = 0;
        pixel_data[90][48] = 0;
        pixel_data[90][49] = 0;
        pixel_data[90][50] = 0;
        pixel_data[90][51] = 0;
        pixel_data[90][52] = 0;
        pixel_data[90][53] = 0;
        pixel_data[90][54] = 0;
        pixel_data[90][55] = 0;
        pixel_data[90][56] = 0;
        pixel_data[90][57] = 0;
        pixel_data[90][58] = 0;
        pixel_data[90][59] = 0;
        pixel_data[90][60] = 0;
        pixel_data[90][61] = 0;
        pixel_data[90][62] = 0;
        pixel_data[90][63] = 0;
        pixel_data[90][64] = 0;
        pixel_data[90][65] = 0;
        pixel_data[90][66] = 0;
        pixel_data[90][67] = 0;
        pixel_data[90][68] = 0;
        pixel_data[90][69] = 0;
        pixel_data[90][70] = 0;
        pixel_data[90][71] = 0;
        pixel_data[90][72] = 0;
        pixel_data[90][73] = 0;
        pixel_data[90][74] = 0;
        pixel_data[90][75] = 0;
        pixel_data[90][76] = 0;
        pixel_data[90][77] = 0;
        pixel_data[90][78] = 0;
        pixel_data[90][79] = 0;
        pixel_data[90][80] = 0;
        pixel_data[90][81] = 0;
        pixel_data[90][82] = 0;
        pixel_data[90][83] = 0;
        pixel_data[90][84] = 0;
        pixel_data[90][85] = 0;
        pixel_data[90][86] = 0;
        pixel_data[90][87] = 0;
        pixel_data[90][88] = 0;
        pixel_data[90][89] = 0;
        pixel_data[90][90] = 0;
        pixel_data[90][91] = 0;
        pixel_data[90][92] = 0;
        pixel_data[90][93] = 0;
        pixel_data[90][94] = 0;
        pixel_data[90][95] = 0;
        pixel_data[90][96] = 0;
        pixel_data[90][97] = 0;
        pixel_data[90][98] = 0;
        pixel_data[90][99] = 0; // y=90
        pixel_data[91][0] = 0;
        pixel_data[91][1] = 0;
        pixel_data[91][2] = 0;
        pixel_data[91][3] = 0;
        pixel_data[91][4] = 0;
        pixel_data[91][5] = 0;
        pixel_data[91][6] = 0;
        pixel_data[91][7] = 0;
        pixel_data[91][8] = 0;
        pixel_data[91][9] = 0;
        pixel_data[91][10] = 0;
        pixel_data[91][11] = 0;
        pixel_data[91][12] = 0;
        pixel_data[91][13] = 0;
        pixel_data[91][14] = 0;
        pixel_data[91][15] = 0;
        pixel_data[91][16] = 0;
        pixel_data[91][17] = 0;
        pixel_data[91][18] = 0;
        pixel_data[91][19] = 0;
        pixel_data[91][20] = 0;
        pixel_data[91][21] = 0;
        pixel_data[91][22] = 0;
        pixel_data[91][23] = 0;
        pixel_data[91][24] = 0;
        pixel_data[91][25] = 0;
        pixel_data[91][26] = 0;
        pixel_data[91][27] = 0;
        pixel_data[91][28] = 0;
        pixel_data[91][29] = 0;
        pixel_data[91][30] = 0;
        pixel_data[91][31] = 0;
        pixel_data[91][32] = 0;
        pixel_data[91][33] = 0;
        pixel_data[91][34] = 0;
        pixel_data[91][35] = 0;
        pixel_data[91][36] = 0;
        pixel_data[91][37] = 0;
        pixel_data[91][38] = 0;
        pixel_data[91][39] = 0;
        pixel_data[91][40] = 0;
        pixel_data[91][41] = 0;
        pixel_data[91][42] = 0;
        pixel_data[91][43] = 0;
        pixel_data[91][44] = 0;
        pixel_data[91][45] = 0;
        pixel_data[91][46] = 0;
        pixel_data[91][47] = 0;
        pixel_data[91][48] = 0;
        pixel_data[91][49] = 0;
        pixel_data[91][50] = 0;
        pixel_data[91][51] = 0;
        pixel_data[91][52] = 0;
        pixel_data[91][53] = 0;
        pixel_data[91][54] = 0;
        pixel_data[91][55] = 0;
        pixel_data[91][56] = 0;
        pixel_data[91][57] = 0;
        pixel_data[91][58] = 0;
        pixel_data[91][59] = 0;
        pixel_data[91][60] = 0;
        pixel_data[91][61] = 0;
        pixel_data[91][62] = 0;
        pixel_data[91][63] = 0;
        pixel_data[91][64] = 0;
        pixel_data[91][65] = 0;
        pixel_data[91][66] = 0;
        pixel_data[91][67] = 0;
        pixel_data[91][68] = 0;
        pixel_data[91][69] = 0;
        pixel_data[91][70] = 0;
        pixel_data[91][71] = 0;
        pixel_data[91][72] = 0;
        pixel_data[91][73] = 0;
        pixel_data[91][74] = 0;
        pixel_data[91][75] = 0;
        pixel_data[91][76] = 0;
        pixel_data[91][77] = 0;
        pixel_data[91][78] = 0;
        pixel_data[91][79] = 0;
        pixel_data[91][80] = 0;
        pixel_data[91][81] = 0;
        pixel_data[91][82] = 0;
        pixel_data[91][83] = 0;
        pixel_data[91][84] = 0;
        pixel_data[91][85] = 0;
        pixel_data[91][86] = 0;
        pixel_data[91][87] = 0;
        pixel_data[91][88] = 0;
        pixel_data[91][89] = 0;
        pixel_data[91][90] = 0;
        pixel_data[91][91] = 0;
        pixel_data[91][92] = 0;
        pixel_data[91][93] = 0;
        pixel_data[91][94] = 0;
        pixel_data[91][95] = 0;
        pixel_data[91][96] = 0;
        pixel_data[91][97] = 0;
        pixel_data[91][98] = 0;
        pixel_data[91][99] = 0; // y=91
        pixel_data[92][0] = 0;
        pixel_data[92][1] = 0;
        pixel_data[92][2] = 0;
        pixel_data[92][3] = 0;
        pixel_data[92][4] = 0;
        pixel_data[92][5] = 0;
        pixel_data[92][6] = 0;
        pixel_data[92][7] = 0;
        pixel_data[92][8] = 0;
        pixel_data[92][9] = 0;
        pixel_data[92][10] = 0;
        pixel_data[92][11] = 0;
        pixel_data[92][12] = 0;
        pixel_data[92][13] = 0;
        pixel_data[92][14] = 0;
        pixel_data[92][15] = 0;
        pixel_data[92][16] = 0;
        pixel_data[92][17] = 0;
        pixel_data[92][18] = 0;
        pixel_data[92][19] = 0;
        pixel_data[92][20] = 0;
        pixel_data[92][21] = 0;
        pixel_data[92][22] = 0;
        pixel_data[92][23] = 0;
        pixel_data[92][24] = 0;
        pixel_data[92][25] = 0;
        pixel_data[92][26] = 0;
        pixel_data[92][27] = 0;
        pixel_data[92][28] = 0;
        pixel_data[92][29] = 0;
        pixel_data[92][30] = 0;
        pixel_data[92][31] = 0;
        pixel_data[92][32] = 0;
        pixel_data[92][33] = 0;
        pixel_data[92][34] = 0;
        pixel_data[92][35] = 0;
        pixel_data[92][36] = 0;
        pixel_data[92][37] = 0;
        pixel_data[92][38] = 0;
        pixel_data[92][39] = 0;
        pixel_data[92][40] = 0;
        pixel_data[92][41] = 0;
        pixel_data[92][42] = 0;
        pixel_data[92][43] = 0;
        pixel_data[92][44] = 0;
        pixel_data[92][45] = 0;
        pixel_data[92][46] = 0;
        pixel_data[92][47] = 0;
        pixel_data[92][48] = 0;
        pixel_data[92][49] = 0;
        pixel_data[92][50] = 0;
        pixel_data[92][51] = 0;
        pixel_data[92][52] = 0;
        pixel_data[92][53] = 0;
        pixel_data[92][54] = 0;
        pixel_data[92][55] = 0;
        pixel_data[92][56] = 0;
        pixel_data[92][57] = 0;
        pixel_data[92][58] = 0;
        pixel_data[92][59] = 0;
        pixel_data[92][60] = 0;
        pixel_data[92][61] = 0;
        pixel_data[92][62] = 0;
        pixel_data[92][63] = 0;
        pixel_data[92][64] = 0;
        pixel_data[92][65] = 0;
        pixel_data[92][66] = 0;
        pixel_data[92][67] = 0;
        pixel_data[92][68] = 0;
        pixel_data[92][69] = 0;
        pixel_data[92][70] = 0;
        pixel_data[92][71] = 0;
        pixel_data[92][72] = 0;
        pixel_data[92][73] = 0;
        pixel_data[92][74] = 0;
        pixel_data[92][75] = 0;
        pixel_data[92][76] = 0;
        pixel_data[92][77] = 0;
        pixel_data[92][78] = 0;
        pixel_data[92][79] = 0;
        pixel_data[92][80] = 0;
        pixel_data[92][81] = 0;
        pixel_data[92][82] = 0;
        pixel_data[92][83] = 0;
        pixel_data[92][84] = 0;
        pixel_data[92][85] = 0;
        pixel_data[92][86] = 0;
        pixel_data[92][87] = 0;
        pixel_data[92][88] = 0;
        pixel_data[92][89] = 0;
        pixel_data[92][90] = 0;
        pixel_data[92][91] = 0;
        pixel_data[92][92] = 0;
        pixel_data[92][93] = 0;
        pixel_data[92][94] = 0;
        pixel_data[92][95] = 0;
        pixel_data[92][96] = 0;
        pixel_data[92][97] = 0;
        pixel_data[92][98] = 0;
        pixel_data[92][99] = 0; // y=92
        pixel_data[93][0] = 0;
        pixel_data[93][1] = 0;
        pixel_data[93][2] = 0;
        pixel_data[93][3] = 0;
        pixel_data[93][4] = 0;
        pixel_data[93][5] = 0;
        pixel_data[93][6] = 0;
        pixel_data[93][7] = 0;
        pixel_data[93][8] = 0;
        pixel_data[93][9] = 0;
        pixel_data[93][10] = 0;
        pixel_data[93][11] = 0;
        pixel_data[93][12] = 0;
        pixel_data[93][13] = 0;
        pixel_data[93][14] = 0;
        pixel_data[93][15] = 0;
        pixel_data[93][16] = 0;
        pixel_data[93][17] = 0;
        pixel_data[93][18] = 0;
        pixel_data[93][19] = 0;
        pixel_data[93][20] = 0;
        pixel_data[93][21] = 0;
        pixel_data[93][22] = 0;
        pixel_data[93][23] = 0;
        pixel_data[93][24] = 0;
        pixel_data[93][25] = 0;
        pixel_data[93][26] = 0;
        pixel_data[93][27] = 0;
        pixel_data[93][28] = 0;
        pixel_data[93][29] = 0;
        pixel_data[93][30] = 0;
        pixel_data[93][31] = 0;
        pixel_data[93][32] = 0;
        pixel_data[93][33] = 0;
        pixel_data[93][34] = 0;
        pixel_data[93][35] = 0;
        pixel_data[93][36] = 0;
        pixel_data[93][37] = 0;
        pixel_data[93][38] = 0;
        pixel_data[93][39] = 0;
        pixel_data[93][40] = 0;
        pixel_data[93][41] = 0;
        pixel_data[93][42] = 0;
        pixel_data[93][43] = 0;
        pixel_data[93][44] = 0;
        pixel_data[93][45] = 0;
        pixel_data[93][46] = 0;
        pixel_data[93][47] = 0;
        pixel_data[93][48] = 0;
        pixel_data[93][49] = 0;
        pixel_data[93][50] = 0;
        pixel_data[93][51] = 0;
        pixel_data[93][52] = 0;
        pixel_data[93][53] = 0;
        pixel_data[93][54] = 0;
        pixel_data[93][55] = 0;
        pixel_data[93][56] = 0;
        pixel_data[93][57] = 0;
        pixel_data[93][58] = 0;
        pixel_data[93][59] = 0;
        pixel_data[93][60] = 0;
        pixel_data[93][61] = 0;
        pixel_data[93][62] = 0;
        pixel_data[93][63] = 0;
        pixel_data[93][64] = 0;
        pixel_data[93][65] = 0;
        pixel_data[93][66] = 0;
        pixel_data[93][67] = 0;
        pixel_data[93][68] = 0;
        pixel_data[93][69] = 0;
        pixel_data[93][70] = 0;
        pixel_data[93][71] = 0;
        pixel_data[93][72] = 0;
        pixel_data[93][73] = 0;
        pixel_data[93][74] = 0;
        pixel_data[93][75] = 0;
        pixel_data[93][76] = 0;
        pixel_data[93][77] = 0;
        pixel_data[93][78] = 0;
        pixel_data[93][79] = 0;
        pixel_data[93][80] = 0;
        pixel_data[93][81] = 0;
        pixel_data[93][82] = 0;
        pixel_data[93][83] = 0;
        pixel_data[93][84] = 0;
        pixel_data[93][85] = 0;
        pixel_data[93][86] = 0;
        pixel_data[93][87] = 0;
        pixel_data[93][88] = 0;
        pixel_data[93][89] = 0;
        pixel_data[93][90] = 0;
        pixel_data[93][91] = 0;
        pixel_data[93][92] = 0;
        pixel_data[93][93] = 0;
        pixel_data[93][94] = 0;
        pixel_data[93][95] = 0;
        pixel_data[93][96] = 0;
        pixel_data[93][97] = 0;
        pixel_data[93][98] = 0;
        pixel_data[93][99] = 0; // y=93
        pixel_data[94][0] = 0;
        pixel_data[94][1] = 0;
        pixel_data[94][2] = 0;
        pixel_data[94][3] = 0;
        pixel_data[94][4] = 0;
        pixel_data[94][5] = 0;
        pixel_data[94][6] = 0;
        pixel_data[94][7] = 0;
        pixel_data[94][8] = 0;
        pixel_data[94][9] = 0;
        pixel_data[94][10] = 0;
        pixel_data[94][11] = 0;
        pixel_data[94][12] = 0;
        pixel_data[94][13] = 0;
        pixel_data[94][14] = 0;
        pixel_data[94][15] = 0;
        pixel_data[94][16] = 0;
        pixel_data[94][17] = 0;
        pixel_data[94][18] = 0;
        pixel_data[94][19] = 0;
        pixel_data[94][20] = 0;
        pixel_data[94][21] = 0;
        pixel_data[94][22] = 0;
        pixel_data[94][23] = 0;
        pixel_data[94][24] = 0;
        pixel_data[94][25] = 0;
        pixel_data[94][26] = 0;
        pixel_data[94][27] = 0;
        pixel_data[94][28] = 0;
        pixel_data[94][29] = 0;
        pixel_data[94][30] = 0;
        pixel_data[94][31] = 0;
        pixel_data[94][32] = 0;
        pixel_data[94][33] = 0;
        pixel_data[94][34] = 0;
        pixel_data[94][35] = 0;
        pixel_data[94][36] = 0;
        pixel_data[94][37] = 0;
        pixel_data[94][38] = 0;
        pixel_data[94][39] = 0;
        pixel_data[94][40] = 0;
        pixel_data[94][41] = 0;
        pixel_data[94][42] = 0;
        pixel_data[94][43] = 0;
        pixel_data[94][44] = 0;
        pixel_data[94][45] = 0;
        pixel_data[94][46] = 0;
        pixel_data[94][47] = 0;
        pixel_data[94][48] = 0;
        pixel_data[94][49] = 0;
        pixel_data[94][50] = 0;
        pixel_data[94][51] = 0;
        pixel_data[94][52] = 0;
        pixel_data[94][53] = 0;
        pixel_data[94][54] = 0;
        pixel_data[94][55] = 0;
        pixel_data[94][56] = 0;
        pixel_data[94][57] = 0;
        pixel_data[94][58] = 0;
        pixel_data[94][59] = 0;
        pixel_data[94][60] = 0;
        pixel_data[94][61] = 0;
        pixel_data[94][62] = 0;
        pixel_data[94][63] = 0;
        pixel_data[94][64] = 0;
        pixel_data[94][65] = 0;
        pixel_data[94][66] = 0;
        pixel_data[94][67] = 0;
        pixel_data[94][68] = 0;
        pixel_data[94][69] = 0;
        pixel_data[94][70] = 0;
        pixel_data[94][71] = 0;
        pixel_data[94][72] = 0;
        pixel_data[94][73] = 0;
        pixel_data[94][74] = 0;
        pixel_data[94][75] = 0;
        pixel_data[94][76] = 0;
        pixel_data[94][77] = 0;
        pixel_data[94][78] = 0;
        pixel_data[94][79] = 0;
        pixel_data[94][80] = 0;
        pixel_data[94][81] = 0;
        pixel_data[94][82] = 0;
        pixel_data[94][83] = 0;
        pixel_data[94][84] = 0;
        pixel_data[94][85] = 0;
        pixel_data[94][86] = 0;
        pixel_data[94][87] = 0;
        pixel_data[94][88] = 0;
        pixel_data[94][89] = 0;
        pixel_data[94][90] = 0;
        pixel_data[94][91] = 0;
        pixel_data[94][92] = 0;
        pixel_data[94][93] = 0;
        pixel_data[94][94] = 0;
        pixel_data[94][95] = 0;
        pixel_data[94][96] = 0;
        pixel_data[94][97] = 0;
        pixel_data[94][98] = 0;
        pixel_data[94][99] = 0; // y=94
        pixel_data[95][0] = 0;
        pixel_data[95][1] = 0;
        pixel_data[95][2] = 0;
        pixel_data[95][3] = 0;
        pixel_data[95][4] = 0;
        pixel_data[95][5] = 0;
        pixel_data[95][6] = 0;
        pixel_data[95][7] = 0;
        pixel_data[95][8] = 0;
        pixel_data[95][9] = 0;
        pixel_data[95][10] = 0;
        pixel_data[95][11] = 0;
        pixel_data[95][12] = 0;
        pixel_data[95][13] = 0;
        pixel_data[95][14] = 0;
        pixel_data[95][15] = 0;
        pixel_data[95][16] = 0;
        pixel_data[95][17] = 0;
        pixel_data[95][18] = 0;
        pixel_data[95][19] = 0;
        pixel_data[95][20] = 0;
        pixel_data[95][21] = 0;
        pixel_data[95][22] = 0;
        pixel_data[95][23] = 0;
        pixel_data[95][24] = 0;
        pixel_data[95][25] = 0;
        pixel_data[95][26] = 0;
        pixel_data[95][27] = 0;
        pixel_data[95][28] = 0;
        pixel_data[95][29] = 0;
        pixel_data[95][30] = 0;
        pixel_data[95][31] = 0;
        pixel_data[95][32] = 0;
        pixel_data[95][33] = 0;
        pixel_data[95][34] = 0;
        pixel_data[95][35] = 0;
        pixel_data[95][36] = 0;
        pixel_data[95][37] = 0;
        pixel_data[95][38] = 0;
        pixel_data[95][39] = 0;
        pixel_data[95][40] = 0;
        pixel_data[95][41] = 0;
        pixel_data[95][42] = 0;
        pixel_data[95][43] = 0;
        pixel_data[95][44] = 0;
        pixel_data[95][45] = 0;
        pixel_data[95][46] = 0;
        pixel_data[95][47] = 0;
        pixel_data[95][48] = 0;
        pixel_data[95][49] = 0;
        pixel_data[95][50] = 0;
        pixel_data[95][51] = 0;
        pixel_data[95][52] = 0;
        pixel_data[95][53] = 0;
        pixel_data[95][54] = 0;
        pixel_data[95][55] = 0;
        pixel_data[95][56] = 0;
        pixel_data[95][57] = 0;
        pixel_data[95][58] = 0;
        pixel_data[95][59] = 0;
        pixel_data[95][60] = 0;
        pixel_data[95][61] = 0;
        pixel_data[95][62] = 0;
        pixel_data[95][63] = 0;
        pixel_data[95][64] = 0;
        pixel_data[95][65] = 0;
        pixel_data[95][66] = 0;
        pixel_data[95][67] = 0;
        pixel_data[95][68] = 0;
        pixel_data[95][69] = 0;
        pixel_data[95][70] = 0;
        pixel_data[95][71] = 0;
        pixel_data[95][72] = 0;
        pixel_data[95][73] = 0;
        pixel_data[95][74] = 0;
        pixel_data[95][75] = 0;
        pixel_data[95][76] = 0;
        pixel_data[95][77] = 0;
        pixel_data[95][78] = 0;
        pixel_data[95][79] = 0;
        pixel_data[95][80] = 0;
        pixel_data[95][81] = 0;
        pixel_data[95][82] = 0;
        pixel_data[95][83] = 0;
        pixel_data[95][84] = 0;
        pixel_data[95][85] = 0;
        pixel_data[95][86] = 0;
        pixel_data[95][87] = 0;
        pixel_data[95][88] = 0;
        pixel_data[95][89] = 0;
        pixel_data[95][90] = 0;
        pixel_data[95][91] = 0;
        pixel_data[95][92] = 0;
        pixel_data[95][93] = 0;
        pixel_data[95][94] = 0;
        pixel_data[95][95] = 0;
        pixel_data[95][96] = 0;
        pixel_data[95][97] = 0;
        pixel_data[95][98] = 0;
        pixel_data[95][99] = 0; // y=95
        pixel_data[96][0] = 0;
        pixel_data[96][1] = 0;
        pixel_data[96][2] = 0;
        pixel_data[96][3] = 0;
        pixel_data[96][4] = 0;
        pixel_data[96][5] = 0;
        pixel_data[96][6] = 0;
        pixel_data[96][7] = 0;
        pixel_data[96][8] = 0;
        pixel_data[96][9] = 0;
        pixel_data[96][10] = 0;
        pixel_data[96][11] = 0;
        pixel_data[96][12] = 0;
        pixel_data[96][13] = 0;
        pixel_data[96][14] = 0;
        pixel_data[96][15] = 0;
        pixel_data[96][16] = 0;
        pixel_data[96][17] = 0;
        pixel_data[96][18] = 0;
        pixel_data[96][19] = 0;
        pixel_data[96][20] = 0;
        pixel_data[96][21] = 0;
        pixel_data[96][22] = 0;
        pixel_data[96][23] = 0;
        pixel_data[96][24] = 0;
        pixel_data[96][25] = 0;
        pixel_data[96][26] = 0;
        pixel_data[96][27] = 0;
        pixel_data[96][28] = 0;
        pixel_data[96][29] = 0;
        pixel_data[96][30] = 0;
        pixel_data[96][31] = 0;
        pixel_data[96][32] = 0;
        pixel_data[96][33] = 0;
        pixel_data[96][34] = 0;
        pixel_data[96][35] = 0;
        pixel_data[96][36] = 0;
        pixel_data[96][37] = 0;
        pixel_data[96][38] = 0;
        pixel_data[96][39] = 0;
        pixel_data[96][40] = 0;
        pixel_data[96][41] = 0;
        pixel_data[96][42] = 0;
        pixel_data[96][43] = 0;
        pixel_data[96][44] = 0;
        pixel_data[96][45] = 0;
        pixel_data[96][46] = 0;
        pixel_data[96][47] = 0;
        pixel_data[96][48] = 0;
        pixel_data[96][49] = 0;
        pixel_data[96][50] = 0;
        pixel_data[96][51] = 0;
        pixel_data[96][52] = 0;
        pixel_data[96][53] = 0;
        pixel_data[96][54] = 0;
        pixel_data[96][55] = 0;
        pixel_data[96][56] = 0;
        pixel_data[96][57] = 0;
        pixel_data[96][58] = 0;
        pixel_data[96][59] = 0;
        pixel_data[96][60] = 0;
        pixel_data[96][61] = 0;
        pixel_data[96][62] = 0;
        pixel_data[96][63] = 0;
        pixel_data[96][64] = 0;
        pixel_data[96][65] = 0;
        pixel_data[96][66] = 0;
        pixel_data[96][67] = 0;
        pixel_data[96][68] = 0;
        pixel_data[96][69] = 0;
        pixel_data[96][70] = 0;
        pixel_data[96][71] = 0;
        pixel_data[96][72] = 0;
        pixel_data[96][73] = 0;
        pixel_data[96][74] = 0;
        pixel_data[96][75] = 0;
        pixel_data[96][76] = 0;
        pixel_data[96][77] = 0;
        pixel_data[96][78] = 0;
        pixel_data[96][79] = 0;
        pixel_data[96][80] = 0;
        pixel_data[96][81] = 0;
        pixel_data[96][82] = 0;
        pixel_data[96][83] = 0;
        pixel_data[96][84] = 0;
        pixel_data[96][85] = 0;
        pixel_data[96][86] = 0;
        pixel_data[96][87] = 0;
        pixel_data[96][88] = 0;
        pixel_data[96][89] = 0;
        pixel_data[96][90] = 0;
        pixel_data[96][91] = 0;
        pixel_data[96][92] = 0;
        pixel_data[96][93] = 0;
        pixel_data[96][94] = 0;
        pixel_data[96][95] = 0;
        pixel_data[96][96] = 0;
        pixel_data[96][97] = 0;
        pixel_data[96][98] = 0;
        pixel_data[96][99] = 0; // y=96
        pixel_data[97][0] = 0;
        pixel_data[97][1] = 0;
        pixel_data[97][2] = 0;
        pixel_data[97][3] = 0;
        pixel_data[97][4] = 0;
        pixel_data[97][5] = 0;
        pixel_data[97][6] = 0;
        pixel_data[97][7] = 0;
        pixel_data[97][8] = 0;
        pixel_data[97][9] = 0;
        pixel_data[97][10] = 0;
        pixel_data[97][11] = 0;
        pixel_data[97][12] = 0;
        pixel_data[97][13] = 0;
        pixel_data[97][14] = 0;
        pixel_data[97][15] = 0;
        pixel_data[97][16] = 0;
        pixel_data[97][17] = 0;
        pixel_data[97][18] = 0;
        pixel_data[97][19] = 0;
        pixel_data[97][20] = 0;
        pixel_data[97][21] = 0;
        pixel_data[97][22] = 0;
        pixel_data[97][23] = 0;
        pixel_data[97][24] = 0;
        pixel_data[97][25] = 0;
        pixel_data[97][26] = 0;
        pixel_data[97][27] = 0;
        pixel_data[97][28] = 0;
        pixel_data[97][29] = 0;
        pixel_data[97][30] = 0;
        pixel_data[97][31] = 0;
        pixel_data[97][32] = 0;
        pixel_data[97][33] = 0;
        pixel_data[97][34] = 0;
        pixel_data[97][35] = 0;
        pixel_data[97][36] = 0;
        pixel_data[97][37] = 0;
        pixel_data[97][38] = 0;
        pixel_data[97][39] = 0;
        pixel_data[97][40] = 0;
        pixel_data[97][41] = 0;
        pixel_data[97][42] = 0;
        pixel_data[97][43] = 0;
        pixel_data[97][44] = 0;
        pixel_data[97][45] = 0;
        pixel_data[97][46] = 0;
        pixel_data[97][47] = 0;
        pixel_data[97][48] = 0;
        pixel_data[97][49] = 0;
        pixel_data[97][50] = 0;
        pixel_data[97][51] = 0;
        pixel_data[97][52] = 0;
        pixel_data[97][53] = 0;
        pixel_data[97][54] = 0;
        pixel_data[97][55] = 0;
        pixel_data[97][56] = 0;
        pixel_data[97][57] = 0;
        pixel_data[97][58] = 0;
        pixel_data[97][59] = 0;
        pixel_data[97][60] = 0;
        pixel_data[97][61] = 0;
        pixel_data[97][62] = 0;
        pixel_data[97][63] = 0;
        pixel_data[97][64] = 0;
        pixel_data[97][65] = 0;
        pixel_data[97][66] = 0;
        pixel_data[97][67] = 0;
        pixel_data[97][68] = 0;
        pixel_data[97][69] = 0;
        pixel_data[97][70] = 0;
        pixel_data[97][71] = 0;
        pixel_data[97][72] = 0;
        pixel_data[97][73] = 0;
        pixel_data[97][74] = 0;
        pixel_data[97][75] = 0;
        pixel_data[97][76] = 0;
        pixel_data[97][77] = 0;
        pixel_data[97][78] = 0;
        pixel_data[97][79] = 0;
        pixel_data[97][80] = 0;
        pixel_data[97][81] = 0;
        pixel_data[97][82] = 0;
        pixel_data[97][83] = 0;
        pixel_data[97][84] = 0;
        pixel_data[97][85] = 0;
        pixel_data[97][86] = 0;
        pixel_data[97][87] = 0;
        pixel_data[97][88] = 0;
        pixel_data[97][89] = 0;
        pixel_data[97][90] = 0;
        pixel_data[97][91] = 0;
        pixel_data[97][92] = 0;
        pixel_data[97][93] = 0;
        pixel_data[97][94] = 0;
        pixel_data[97][95] = 0;
        pixel_data[97][96] = 0;
        pixel_data[97][97] = 0;
        pixel_data[97][98] = 0;
        pixel_data[97][99] = 0; // y=97
        pixel_data[98][0] = 0;
        pixel_data[98][1] = 0;
        pixel_data[98][2] = 0;
        pixel_data[98][3] = 0;
        pixel_data[98][4] = 0;
        pixel_data[98][5] = 0;
        pixel_data[98][6] = 0;
        pixel_data[98][7] = 0;
        pixel_data[98][8] = 0;
        pixel_data[98][9] = 0;
        pixel_data[98][10] = 0;
        pixel_data[98][11] = 0;
        pixel_data[98][12] = 0;
        pixel_data[98][13] = 0;
        pixel_data[98][14] = 0;
        pixel_data[98][15] = 0;
        pixel_data[98][16] = 0;
        pixel_data[98][17] = 0;
        pixel_data[98][18] = 0;
        pixel_data[98][19] = 0;
        pixel_data[98][20] = 0;
        pixel_data[98][21] = 0;
        pixel_data[98][22] = 0;
        pixel_data[98][23] = 0;
        pixel_data[98][24] = 0;
        pixel_data[98][25] = 0;
        pixel_data[98][26] = 0;
        pixel_data[98][27] = 0;
        pixel_data[98][28] = 0;
        pixel_data[98][29] = 0;
        pixel_data[98][30] = 0;
        pixel_data[98][31] = 0;
        pixel_data[98][32] = 0;
        pixel_data[98][33] = 0;
        pixel_data[98][34] = 0;
        pixel_data[98][35] = 0;
        pixel_data[98][36] = 0;
        pixel_data[98][37] = 0;
        pixel_data[98][38] = 0;
        pixel_data[98][39] = 0;
        pixel_data[98][40] = 0;
        pixel_data[98][41] = 0;
        pixel_data[98][42] = 0;
        pixel_data[98][43] = 0;
        pixel_data[98][44] = 0;
        pixel_data[98][45] = 0;
        pixel_data[98][46] = 0;
        pixel_data[98][47] = 0;
        pixel_data[98][48] = 0;
        pixel_data[98][49] = 0;
        pixel_data[98][50] = 0;
        pixel_data[98][51] = 0;
        pixel_data[98][52] = 0;
        pixel_data[98][53] = 0;
        pixel_data[98][54] = 0;
        pixel_data[98][55] = 0;
        pixel_data[98][56] = 0;
        pixel_data[98][57] = 0;
        pixel_data[98][58] = 0;
        pixel_data[98][59] = 0;
        pixel_data[98][60] = 0;
        pixel_data[98][61] = 0;
        pixel_data[98][62] = 0;
        pixel_data[98][63] = 0;
        pixel_data[98][64] = 0;
        pixel_data[98][65] = 0;
        pixel_data[98][66] = 0;
        pixel_data[98][67] = 0;
        pixel_data[98][68] = 0;
        pixel_data[98][69] = 0;
        pixel_data[98][70] = 0;
        pixel_data[98][71] = 0;
        pixel_data[98][72] = 0;
        pixel_data[98][73] = 0;
        pixel_data[98][74] = 0;
        pixel_data[98][75] = 0;
        pixel_data[98][76] = 0;
        pixel_data[98][77] = 0;
        pixel_data[98][78] = 0;
        pixel_data[98][79] = 0;
        pixel_data[98][80] = 0;
        pixel_data[98][81] = 0;
        pixel_data[98][82] = 0;
        pixel_data[98][83] = 0;
        pixel_data[98][84] = 0;
        pixel_data[98][85] = 0;
        pixel_data[98][86] = 0;
        pixel_data[98][87] = 0;
        pixel_data[98][88] = 0;
        pixel_data[98][89] = 0;
        pixel_data[98][90] = 0;
        pixel_data[98][91] = 0;
        pixel_data[98][92] = 0;
        pixel_data[98][93] = 0;
        pixel_data[98][94] = 0;
        pixel_data[98][95] = 0;
        pixel_data[98][96] = 0;
        pixel_data[98][97] = 0;
        pixel_data[98][98] = 0;
        pixel_data[98][99] = 0; // y=98
        pixel_data[99][0] = 0;
        pixel_data[99][1] = 0;
        pixel_data[99][2] = 0;
        pixel_data[99][3] = 0;
        pixel_data[99][4] = 0;
        pixel_data[99][5] = 0;
        pixel_data[99][6] = 0;
        pixel_data[99][7] = 0;
        pixel_data[99][8] = 0;
        pixel_data[99][9] = 0;
        pixel_data[99][10] = 0;
        pixel_data[99][11] = 0;
        pixel_data[99][12] = 0;
        pixel_data[99][13] = 0;
        pixel_data[99][14] = 0;
        pixel_data[99][15] = 0;
        pixel_data[99][16] = 0;
        pixel_data[99][17] = 0;
        pixel_data[99][18] = 0;
        pixel_data[99][19] = 0;
        pixel_data[99][20] = 0;
        pixel_data[99][21] = 0;
        pixel_data[99][22] = 0;
        pixel_data[99][23] = 0;
        pixel_data[99][24] = 0;
        pixel_data[99][25] = 0;
        pixel_data[99][26] = 0;
        pixel_data[99][27] = 0;
        pixel_data[99][28] = 0;
        pixel_data[99][29] = 0;
        pixel_data[99][30] = 0;
        pixel_data[99][31] = 0;
        pixel_data[99][32] = 0;
        pixel_data[99][33] = 0;
        pixel_data[99][34] = 0;
        pixel_data[99][35] = 0;
        pixel_data[99][36] = 0;
        pixel_data[99][37] = 0;
        pixel_data[99][38] = 0;
        pixel_data[99][39] = 0;
        pixel_data[99][40] = 0;
        pixel_data[99][41] = 0;
        pixel_data[99][42] = 0;
        pixel_data[99][43] = 0;
        pixel_data[99][44] = 0;
        pixel_data[99][45] = 0;
        pixel_data[99][46] = 0;
        pixel_data[99][47] = 0;
        pixel_data[99][48] = 0;
        pixel_data[99][49] = 0;
        pixel_data[99][50] = 0;
        pixel_data[99][51] = 0;
        pixel_data[99][52] = 0;
        pixel_data[99][53] = 0;
        pixel_data[99][54] = 0;
        pixel_data[99][55] = 0;
        pixel_data[99][56] = 0;
        pixel_data[99][57] = 0;
        pixel_data[99][58] = 0;
        pixel_data[99][59] = 0;
        pixel_data[99][60] = 0;
        pixel_data[99][61] = 0;
        pixel_data[99][62] = 0;
        pixel_data[99][63] = 0;
        pixel_data[99][64] = 0;
        pixel_data[99][65] = 0;
        pixel_data[99][66] = 0;
        pixel_data[99][67] = 0;
        pixel_data[99][68] = 0;
        pixel_data[99][69] = 0;
        pixel_data[99][70] = 0;
        pixel_data[99][71] = 0;
        pixel_data[99][72] = 0;
        pixel_data[99][73] = 0;
        pixel_data[99][74] = 0;
        pixel_data[99][75] = 0;
        pixel_data[99][76] = 0;
        pixel_data[99][77] = 0;
        pixel_data[99][78] = 0;
        pixel_data[99][79] = 0;
        pixel_data[99][80] = 0;
        pixel_data[99][81] = 0;
        pixel_data[99][82] = 0;
        pixel_data[99][83] = 0;
        pixel_data[99][84] = 0;
        pixel_data[99][85] = 0;
        pixel_data[99][86] = 0;
        pixel_data[99][87] = 0;
        pixel_data[99][88] = 0;
        pixel_data[99][89] = 0;
        pixel_data[99][90] = 0;
        pixel_data[99][91] = 0;
        pixel_data[99][92] = 0;
        pixel_data[99][93] = 0;
        pixel_data[99][94] = 0;
        pixel_data[99][95] = 0;
        pixel_data[99][96] = 0;
        pixel_data[99][97] = 0;
        pixel_data[99][98] = 0;
        pixel_data[99][99] = 0; // y=99
    end
endmodule
