module player1_shield_lut(output reg [3:0] pixel_data [0:49][0:49]);
    initial begin
        pixel_data[0][0] = 0;
        pixel_data[0][1] = 0;
        pixel_data[0][2] = 0;
        pixel_data[0][3] = 0;
        pixel_data[0][4] = 0;
        pixel_data[0][5] = 0;
        pixel_data[0][6] = 0;
        pixel_data[0][7] = 0;
        pixel_data[0][8] = 0;
        pixel_data[0][9] = 0;
        pixel_data[0][10] = 0;
        pixel_data[0][11] = 0;
        pixel_data[0][12] = 0;
        pixel_data[0][13] = 0;
        pixel_data[0][14] = 0;
        pixel_data[0][15] = 0;
        pixel_data[0][16] = 0;
        pixel_data[0][17] = 0;
        pixel_data[0][18] = 0;
        pixel_data[0][19] = 2;
        pixel_data[0][20] = 11;
        pixel_data[0][21] = 10;
        pixel_data[0][22] = 10;
        pixel_data[0][23] = 7;
        pixel_data[0][24] = 11;
        pixel_data[0][25] = 11;
        pixel_data[0][26] = 11;
        pixel_data[0][27] = 11;
        pixel_data[0][28] = 11;
        pixel_data[0][29] = 7;
        pixel_data[0][30] = 7;
        pixel_data[0][31] = 5;
        pixel_data[0][32] = 0;
        pixel_data[0][33] = 0;
        pixel_data[0][34] = 0;
        pixel_data[0][35] = 0;
        pixel_data[0][36] = 0;
        pixel_data[0][37] = 0;
        pixel_data[0][38] = 0;
        pixel_data[0][39] = 0;
        pixel_data[0][40] = 0;
        pixel_data[0][41] = 0;
        pixel_data[0][42] = 0;
        pixel_data[0][43] = 0;
        pixel_data[0][44] = 0;
        pixel_data[0][45] = 0;
        pixel_data[0][46] = 0;
        pixel_data[0][47] = 0;
        pixel_data[0][48] = 0;
        pixel_data[0][49] = 0; // y=0
        pixel_data[1][0] = 0;
        pixel_data[1][1] = 0;
        pixel_data[1][2] = 0;
        pixel_data[1][3] = 0;
        pixel_data[1][4] = 0;
        pixel_data[1][5] = 0;
        pixel_data[1][6] = 0;
        pixel_data[1][7] = 0;
        pixel_data[1][8] = 0;
        pixel_data[1][9] = 0;
        pixel_data[1][10] = 0;
        pixel_data[1][11] = 0;
        pixel_data[1][12] = 0;
        pixel_data[1][13] = 0;
        pixel_data[1][14] = 0;
        pixel_data[1][15] = 0;
        pixel_data[1][16] = 2;
        pixel_data[1][17] = 12;
        pixel_data[1][18] = 1;
        pixel_data[1][19] = 0;
        pixel_data[1][20] = 0;
        pixel_data[1][21] = 0;
        pixel_data[1][22] = 0;
        pixel_data[1][23] = 0;
        pixel_data[1][24] = 0;
        pixel_data[1][25] = 0;
        pixel_data[1][26] = 0;
        pixel_data[1][27] = 0;
        pixel_data[1][28] = 0;
        pixel_data[1][29] = 0;
        pixel_data[1][30] = 0;
        pixel_data[1][31] = 0;
        pixel_data[1][32] = 2;
        pixel_data[1][33] = 1;
        pixel_data[1][34] = 5;
        pixel_data[1][35] = 0;
        pixel_data[1][36] = 0;
        pixel_data[1][37] = 0;
        pixel_data[1][38] = 0;
        pixel_data[1][39] = 0;
        pixel_data[1][40] = 0;
        pixel_data[1][41] = 0;
        pixel_data[1][42] = 0;
        pixel_data[1][43] = 0;
        pixel_data[1][44] = 0;
        pixel_data[1][45] = 0;
        pixel_data[1][46] = 0;
        pixel_data[1][47] = 0;
        pixel_data[1][48] = 0;
        pixel_data[1][49] = 0; // y=1
        pixel_data[2][0] = 0;
        pixel_data[2][1] = 0;
        pixel_data[2][2] = 0;
        pixel_data[2][3] = 0;
        pixel_data[2][4] = 0;
        pixel_data[2][5] = 0;
        pixel_data[2][6] = 0;
        pixel_data[2][7] = 0;
        pixel_data[2][8] = 0;
        pixel_data[2][9] = 0;
        pixel_data[2][10] = 0;
        pixel_data[2][11] = 0;
        pixel_data[2][12] = 0;
        pixel_data[2][13] = 0;
        pixel_data[2][14] = 2;
        pixel_data[2][15] = 11;
        pixel_data[2][16] = 0;
        pixel_data[2][17] = 0;
        pixel_data[2][18] = 0;
        pixel_data[2][19] = 2;
        pixel_data[2][20] = 13;
        pixel_data[2][21] = 13;
        pixel_data[2][22] = 11;
        pixel_data[2][23] = 10;
        pixel_data[2][24] = 10;
        pixel_data[2][25] = 10;
        pixel_data[2][26] = 10;
        pixel_data[2][27] = 10;
        pixel_data[2][28] = 15;
        pixel_data[2][29] = 14;
        pixel_data[2][30] = 10;
        pixel_data[2][31] = 14;
        pixel_data[2][32] = 0;
        pixel_data[2][33] = 0;
        pixel_data[2][34] = 0;
        pixel_data[2][35] = 2;
        pixel_data[2][36] = 5;
        pixel_data[2][37] = 0;
        pixel_data[2][38] = 0;
        pixel_data[2][39] = 0;
        pixel_data[2][40] = 0;
        pixel_data[2][41] = 0;
        pixel_data[2][42] = 0;
        pixel_data[2][43] = 0;
        pixel_data[2][44] = 0;
        pixel_data[2][45] = 0;
        pixel_data[2][46] = 0;
        pixel_data[2][47] = 0;
        pixel_data[2][48] = 0;
        pixel_data[2][49] = 0; // y=2
        pixel_data[3][0] = 0;
        pixel_data[3][1] = 0;
        pixel_data[3][2] = 0;
        pixel_data[3][3] = 0;
        pixel_data[3][4] = 0;
        pixel_data[3][5] = 0;
        pixel_data[3][6] = 0;
        pixel_data[3][7] = 0;
        pixel_data[3][8] = 0;
        pixel_data[3][9] = 0;
        pixel_data[3][10] = 0;
        pixel_data[3][11] = 0;
        pixel_data[3][12] = 0;
        pixel_data[3][13] = 2;
        pixel_data[3][14] = 0;
        pixel_data[3][15] = 0;
        pixel_data[3][16] = 2;
        pixel_data[3][17] = 1;
        pixel_data[3][18] = 11;
        pixel_data[3][19] = 11;
        pixel_data[3][20] = 6;
        pixel_data[3][21] = 4;
        pixel_data[3][22] = 4;
        pixel_data[3][23] = 4;
        pixel_data[3][24] = 4;
        pixel_data[3][25] = 4;
        pixel_data[3][26] = 4;
        pixel_data[3][27] = 6;
        pixel_data[3][28] = 9;
        pixel_data[3][29] = 10;
        pixel_data[3][30] = 10;
        pixel_data[3][31] = 9;
        pixel_data[3][32] = 15;
        pixel_data[3][33] = 14;
        pixel_data[3][34] = 14;
        pixel_data[3][35] = 0;
        pixel_data[3][36] = 0;
        pixel_data[3][37] = 5;
        pixel_data[3][38] = 5;
        pixel_data[3][39] = 0;
        pixel_data[3][40] = 0;
        pixel_data[3][41] = 0;
        pixel_data[3][42] = 0;
        pixel_data[3][43] = 0;
        pixel_data[3][44] = 0;
        pixel_data[3][45] = 0;
        pixel_data[3][46] = 0;
        pixel_data[3][47] = 0;
        pixel_data[3][48] = 0;
        pixel_data[3][49] = 0; // y=3
        pixel_data[4][0] = 0;
        pixel_data[4][1] = 0;
        pixel_data[4][2] = 0;
        pixel_data[4][3] = 0;
        pixel_data[4][4] = 0;
        pixel_data[4][5] = 0;
        pixel_data[4][6] = 0;
        pixel_data[4][7] = 0;
        pixel_data[4][8] = 0;
        pixel_data[4][9] = 0;
        pixel_data[4][10] = 0;
        pixel_data[4][11] = 0;
        pixel_data[4][12] = 10;
        pixel_data[4][13] = 0;
        pixel_data[4][14] = 2;
        pixel_data[4][15] = 11;
        pixel_data[4][16] = 9;
        pixel_data[4][17] = 9;
        pixel_data[4][18] = 3;
        pixel_data[4][19] = 15;
        pixel_data[4][20] = 15;
        pixel_data[4][21] = 15;
        pixel_data[4][22] = 15;
        pixel_data[4][23] = 4;
        pixel_data[4][24] = 3;
        pixel_data[4][25] = 4;
        pixel_data[4][26] = 3;
        pixel_data[4][27] = 3;
        pixel_data[4][28] = 3;
        pixel_data[4][29] = 3;
        pixel_data[4][30] = 15;
        pixel_data[4][31] = 6;
        pixel_data[4][32] = 9;
        pixel_data[4][33] = 6;
        pixel_data[4][34] = 10;
        pixel_data[4][35] = 14;
        pixel_data[4][36] = 14;
        pixel_data[4][37] = 0;
        pixel_data[4][38] = 0;
        pixel_data[4][39] = 5;
        pixel_data[4][40] = 0;
        pixel_data[4][41] = 0;
        pixel_data[4][42] = 0;
        pixel_data[4][43] = 0;
        pixel_data[4][44] = 0;
        pixel_data[4][45] = 0;
        pixel_data[4][46] = 0;
        pixel_data[4][47] = 0;
        pixel_data[4][48] = 0;
        pixel_data[4][49] = 0; // y=4
        pixel_data[5][0] = 0;
        pixel_data[5][1] = 0;
        pixel_data[5][2] = 0;
        pixel_data[5][3] = 0;
        pixel_data[5][4] = 0;
        pixel_data[5][5] = 0;
        pixel_data[5][6] = 0;
        pixel_data[5][7] = 0;
        pixel_data[5][8] = 0;
        pixel_data[5][9] = 0;
        pixel_data[5][10] = 0;
        pixel_data[5][11] = 7;
        pixel_data[5][12] = 0;
        pixel_data[5][13] = 2;
        pixel_data[5][14] = 11;
        pixel_data[5][15] = 6;
        pixel_data[5][16] = 15;
        pixel_data[5][17] = 15;
        pixel_data[5][18] = 15;
        pixel_data[5][19] = 15;
        pixel_data[5][20] = 15;
        pixel_data[5][21] = 15;
        pixel_data[5][22] = 15;
        pixel_data[5][23] = 4;
        pixel_data[5][24] = 4;
        pixel_data[5][25] = 4;
        pixel_data[5][26] = 4;
        pixel_data[5][27] = 4;
        pixel_data[5][28] = 4;
        pixel_data[5][29] = 4;
        pixel_data[5][30] = 4;
        pixel_data[5][31] = 3;
        pixel_data[5][32] = 15;
        pixel_data[5][33] = 15;
        pixel_data[5][34] = 6;
        pixel_data[5][35] = 9;
        pixel_data[5][36] = 9;
        pixel_data[5][37] = 14;
        pixel_data[5][38] = 14;
        pixel_data[5][39] = 0;
        pixel_data[5][40] = 5;
        pixel_data[5][41] = 0;
        pixel_data[5][42] = 0;
        pixel_data[5][43] = 0;
        pixel_data[5][44] = 0;
        pixel_data[5][45] = 0;
        pixel_data[5][46] = 0;
        pixel_data[5][47] = 0;
        pixel_data[5][48] = 0;
        pixel_data[5][49] = 0; // y=5
        pixel_data[6][0] = 0;
        pixel_data[6][1] = 0;
        pixel_data[6][2] = 0;
        pixel_data[6][3] = 0;
        pixel_data[6][4] = 0;
        pixel_data[6][5] = 0;
        pixel_data[6][6] = 0;
        pixel_data[6][7] = 0;
        pixel_data[6][8] = 0;
        pixel_data[6][9] = 2;
        pixel_data[6][10] = 11;
        pixel_data[6][11] = 2;
        pixel_data[6][12] = 13;
        pixel_data[6][13] = 10;
        pixel_data[6][14] = 3;
        pixel_data[6][15] = 15;
        pixel_data[6][16] = 15;
        pixel_data[6][17] = 15;
        pixel_data[6][18] = 15;
        pixel_data[6][19] = 15;
        pixel_data[6][20] = 15;
        pixel_data[6][21] = 15;
        pixel_data[6][22] = 15;
        pixel_data[6][23] = 4;
        pixel_data[6][24] = 4;
        pixel_data[6][25] = 4;
        pixel_data[6][26] = 4;
        pixel_data[6][27] = 4;
        pixel_data[6][28] = 4;
        pixel_data[6][29] = 4;
        pixel_data[6][30] = 4;
        pixel_data[6][31] = 4;
        pixel_data[6][32] = 4;
        pixel_data[6][33] = 4;
        pixel_data[6][34] = 15;
        pixel_data[6][35] = 6;
        pixel_data[6][36] = 9;
        pixel_data[6][37] = 9;
        pixel_data[6][38] = 14;
        pixel_data[6][39] = 14;
        pixel_data[6][40] = 0;
        pixel_data[6][41] = 5;
        pixel_data[6][42] = 0;
        pixel_data[6][43] = 0;
        pixel_data[6][44] = 0;
        pixel_data[6][45] = 0;
        pixel_data[6][46] = 0;
        pixel_data[6][47] = 0;
        pixel_data[6][48] = 0;
        pixel_data[6][49] = 0; // y=6
        pixel_data[7][0] = 0;
        pixel_data[7][1] = 0;
        pixel_data[7][2] = 0;
        pixel_data[7][3] = 0;
        pixel_data[7][4] = 0;
        pixel_data[7][5] = 0;
        pixel_data[7][6] = 0;
        pixel_data[7][7] = 0;
        pixel_data[7][8] = 0;
        pixel_data[7][9] = 12;
        pixel_data[7][10] = 0;
        pixel_data[7][11] = 13;
        pixel_data[7][12] = 9;
        pixel_data[7][13] = 15;
        pixel_data[7][14] = 15;
        pixel_data[7][15] = 15;
        pixel_data[7][16] = 15;
        pixel_data[7][17] = 15;
        pixel_data[7][18] = 15;
        pixel_data[7][19] = 15;
        pixel_data[7][20] = 15;
        pixel_data[7][21] = 5;
        pixel_data[7][22] = 4;
        pixel_data[7][23] = 4;
        pixel_data[7][24] = 4;
        pixel_data[7][25] = 4;
        pixel_data[7][26] = 4;
        pixel_data[7][27] = 4;
        pixel_data[7][28] = 4;
        pixel_data[7][29] = 4;
        pixel_data[7][30] = 4;
        pixel_data[7][31] = 4;
        pixel_data[7][32] = 4;
        pixel_data[7][33] = 4;
        pixel_data[7][34] = 4;
        pixel_data[7][35] = 3;
        pixel_data[7][36] = 3;
        pixel_data[7][37] = 9;
        pixel_data[7][38] = 10;
        pixel_data[7][39] = 14;
        pixel_data[7][40] = 14;
        pixel_data[7][41] = 0;
        pixel_data[7][42] = 5;
        pixel_data[7][43] = 0;
        pixel_data[7][44] = 0;
        pixel_data[7][45] = 0;
        pixel_data[7][46] = 0;
        pixel_data[7][47] = 0;
        pixel_data[7][48] = 0;
        pixel_data[7][49] = 0; // y=7
        pixel_data[8][0] = 0;
        pixel_data[8][1] = 0;
        pixel_data[8][2] = 0;
        pixel_data[8][3] = 0;
        pixel_data[8][4] = 0;
        pixel_data[8][5] = 0;
        pixel_data[8][6] = 0;
        pixel_data[8][7] = 0;
        pixel_data[8][8] = 10;
        pixel_data[8][9] = 0;
        pixel_data[8][10] = 12;
        pixel_data[8][11] = 9;
        pixel_data[8][12] = 15;
        pixel_data[8][13] = 15;
        pixel_data[8][14] = 15;
        pixel_data[8][15] = 15;
        pixel_data[8][16] = 15;
        pixel_data[8][17] = 15;
        pixel_data[8][18] = 15;
        pixel_data[8][19] = 15;
        pixel_data[8][20] = 3;
        pixel_data[8][21] = 4;
        pixel_data[8][22] = 4;
        pixel_data[8][23] = 4;
        pixel_data[8][24] = 4;
        pixel_data[8][25] = 4;
        pixel_data[8][26] = 4;
        pixel_data[8][27] = 4;
        pixel_data[8][28] = 4;
        pixel_data[8][29] = 4;
        pixel_data[8][30] = 4;
        pixel_data[8][31] = 4;
        pixel_data[8][32] = 4;
        pixel_data[8][33] = 4;
        pixel_data[8][34] = 4;
        pixel_data[8][35] = 4;
        pixel_data[8][36] = 4;
        pixel_data[8][37] = 3;
        pixel_data[8][38] = 6;
        pixel_data[8][39] = 10;
        pixel_data[8][40] = 14;
        pixel_data[8][41] = 14;
        pixel_data[8][42] = 0;
        pixel_data[8][43] = 5;
        pixel_data[8][44] = 0;
        pixel_data[8][45] = 0;
        pixel_data[8][46] = 0;
        pixel_data[8][47] = 0;
        pixel_data[8][48] = 0;
        pixel_data[8][49] = 0; // y=8
        pixel_data[9][0] = 0;
        pixel_data[9][1] = 0;
        pixel_data[9][2] = 0;
        pixel_data[9][3] = 0;
        pixel_data[9][4] = 0;
        pixel_data[9][5] = 0;
        pixel_data[9][6] = 0;
        pixel_data[9][7] = 12;
        pixel_data[9][8] = 0;
        pixel_data[9][9] = 12;
        pixel_data[9][10] = 9;
        pixel_data[9][11] = 15;
        pixel_data[9][12] = 15;
        pixel_data[9][13] = 15;
        pixel_data[9][14] = 15;
        pixel_data[9][15] = 15;
        pixel_data[9][16] = 15;
        pixel_data[9][17] = 15;
        pixel_data[9][18] = 15;
        pixel_data[9][19] = 3;
        pixel_data[9][20] = 4;
        pixel_data[9][21] = 4;
        pixel_data[9][22] = 4;
        pixel_data[9][23] = 4;
        pixel_data[9][24] = 4;
        pixel_data[9][25] = 4;
        pixel_data[9][26] = 4;
        pixel_data[9][27] = 4;
        pixel_data[9][28] = 4;
        pixel_data[9][29] = 4;
        pixel_data[9][30] = 4;
        pixel_data[9][31] = 4;
        pixel_data[9][32] = 4;
        pixel_data[9][33] = 4;
        pixel_data[9][34] = 4;
        pixel_data[9][35] = 4;
        pixel_data[9][36] = 4;
        pixel_data[9][37] = 4;
        pixel_data[9][38] = 15;
        pixel_data[9][39] = 6;
        pixel_data[9][40] = 10;
        pixel_data[9][41] = 14;
        pixel_data[9][42] = 14;
        pixel_data[9][43] = 0;
        pixel_data[9][44] = 5;
        pixel_data[9][45] = 0;
        pixel_data[9][46] = 0;
        pixel_data[9][47] = 0;
        pixel_data[9][48] = 0;
        pixel_data[9][49] = 0; // y=9
        pixel_data[10][0] = 0;
        pixel_data[10][1] = 0;
        pixel_data[10][2] = 0;
        pixel_data[10][3] = 0;
        pixel_data[10][4] = 0;
        pixel_data[10][5] = 0;
        pixel_data[10][6] = 11;
        pixel_data[10][7] = 2;
        pixel_data[10][8] = 10;
        pixel_data[10][9] = 9;
        pixel_data[10][10] = 4;
        pixel_data[10][11] = 15;
        pixel_data[10][12] = 15;
        pixel_data[10][13] = 15;
        pixel_data[10][14] = 15;
        pixel_data[10][15] = 15;
        pixel_data[10][16] = 15;
        pixel_data[10][17] = 15;
        pixel_data[10][18] = 3;
        pixel_data[10][19] = 4;
        pixel_data[10][20] = 4;
        pixel_data[10][21] = 4;
        pixel_data[10][22] = 4;
        pixel_data[10][23] = 4;
        pixel_data[10][24] = 4;
        pixel_data[10][25] = 4;
        pixel_data[10][26] = 4;
        pixel_data[10][27] = 4;
        pixel_data[10][28] = 4;
        pixel_data[10][29] = 4;
        pixel_data[10][30] = 4;
        pixel_data[10][31] = 4;
        pixel_data[10][32] = 4;
        pixel_data[10][33] = 4;
        pixel_data[10][34] = 4;
        pixel_data[10][35] = 4;
        pixel_data[10][36] = 4;
        pixel_data[10][37] = 4;
        pixel_data[10][38] = 4;
        pixel_data[10][39] = 3;
        pixel_data[10][40] = 9;
        pixel_data[10][41] = 9;
        pixel_data[10][42] = 14;
        pixel_data[10][43] = 14;
        pixel_data[10][44] = 0;
        pixel_data[10][45] = 5;
        pixel_data[10][46] = 0;
        pixel_data[10][47] = 0;
        pixel_data[10][48] = 0;
        pixel_data[10][49] = 0; // y=10
        pixel_data[11][0] = 0;
        pixel_data[11][1] = 0;
        pixel_data[11][2] = 0;
        pixel_data[11][3] = 0;
        pixel_data[11][4] = 0;
        pixel_data[11][5] = 5;
        pixel_data[11][6] = 11;
        pixel_data[11][7] = 0;
        pixel_data[11][8] = 10;
        pixel_data[11][9] = 6;
        pixel_data[11][10] = 15;
        pixel_data[11][11] = 15;
        pixel_data[11][12] = 15;
        pixel_data[11][13] = 15;
        pixel_data[11][14] = 15;
        pixel_data[11][15] = 15;
        pixel_data[11][16] = 15;
        pixel_data[11][17] = 4;
        pixel_data[11][18] = 4;
        pixel_data[11][19] = 4;
        pixel_data[11][20] = 4;
        pixel_data[11][21] = 4;
        pixel_data[11][22] = 4;
        pixel_data[11][23] = 4;
        pixel_data[11][24] = 4;
        pixel_data[11][25] = 4;
        pixel_data[11][26] = 4;
        pixel_data[11][27] = 4;
        pixel_data[11][28] = 4;
        pixel_data[11][29] = 4;
        pixel_data[11][30] = 4;
        pixel_data[11][31] = 4;
        pixel_data[11][32] = 4;
        pixel_data[11][33] = 4;
        pixel_data[11][34] = 4;
        pixel_data[11][35] = 4;
        pixel_data[11][36] = 4;
        pixel_data[11][37] = 4;
        pixel_data[11][38] = 4;
        pixel_data[11][39] = 4;
        pixel_data[11][40] = 15;
        pixel_data[11][41] = 9;
        pixel_data[11][42] = 14;
        pixel_data[11][43] = 14;
        pixel_data[11][44] = 15;
        pixel_data[11][45] = 0;
        pixel_data[11][46] = 5;
        pixel_data[11][47] = 0;
        pixel_data[11][48] = 0;
        pixel_data[11][49] = 0; // y=11
        pixel_data[12][0] = 0;
        pixel_data[12][1] = 0;
        pixel_data[12][2] = 0;
        pixel_data[12][3] = 0;
        pixel_data[12][4] = 0;
        pixel_data[12][5] = 11;
        pixel_data[12][6] = 0;
        pixel_data[12][7] = 10;
        pixel_data[12][8] = 9;
        pixel_data[12][9] = 15;
        pixel_data[12][10] = 15;
        pixel_data[12][11] = 15;
        pixel_data[12][12] = 15;
        pixel_data[12][13] = 15;
        pixel_data[12][14] = 15;
        pixel_data[12][15] = 15;
        pixel_data[12][16] = 4;
        pixel_data[12][17] = 4;
        pixel_data[12][18] = 4;
        pixel_data[12][19] = 4;
        pixel_data[12][20] = 4;
        pixel_data[12][21] = 4;
        pixel_data[12][22] = 4;
        pixel_data[12][23] = 4;
        pixel_data[12][24] = 4;
        pixel_data[12][25] = 4;
        pixel_data[12][26] = 4;
        pixel_data[12][27] = 4;
        pixel_data[12][28] = 4;
        pixel_data[12][29] = 4;
        pixel_data[12][30] = 4;
        pixel_data[12][31] = 4;
        pixel_data[12][32] = 4;
        pixel_data[12][33] = 4;
        pixel_data[12][34] = 4;
        pixel_data[12][35] = 4;
        pixel_data[12][36] = 4;
        pixel_data[12][37] = 4;
        pixel_data[12][38] = 4;
        pixel_data[12][39] = 4;
        pixel_data[12][40] = 3;
        pixel_data[12][41] = 4;
        pixel_data[12][42] = 9;
        pixel_data[12][43] = 14;
        pixel_data[12][44] = 14;
        pixel_data[12][45] = 2;
        pixel_data[12][46] = 5;
        pixel_data[12][47] = 0;
        pixel_data[12][48] = 0;
        pixel_data[12][49] = 0; // y=12
        pixel_data[13][0] = 0;
        pixel_data[13][1] = 0;
        pixel_data[13][2] = 0;
        pixel_data[13][3] = 0;
        pixel_data[13][4] = 11;
        pixel_data[13][5] = 0;
        pixel_data[13][6] = 10;
        pixel_data[13][7] = 10;
        pixel_data[13][8] = 4;
        pixel_data[13][9] = 15;
        pixel_data[13][10] = 15;
        pixel_data[13][11] = 15;
        pixel_data[13][12] = 15;
        pixel_data[13][13] = 15;
        pixel_data[13][14] = 3;
        pixel_data[13][15] = 4;
        pixel_data[13][16] = 4;
        pixel_data[13][17] = 4;
        pixel_data[13][18] = 4;
        pixel_data[13][19] = 4;
        pixel_data[13][20] = 4;
        pixel_data[13][21] = 4;
        pixel_data[13][22] = 4;
        pixel_data[13][23] = 4;
        pixel_data[13][24] = 4;
        pixel_data[13][25] = 4;
        pixel_data[13][26] = 4;
        pixel_data[13][27] = 4;
        pixel_data[13][28] = 4;
        pixel_data[13][29] = 4;
        pixel_data[13][30] = 4;
        pixel_data[13][31] = 4;
        pixel_data[13][32] = 4;
        pixel_data[13][33] = 4;
        pixel_data[13][34] = 4;
        pixel_data[13][35] = 4;
        pixel_data[13][36] = 4;
        pixel_data[13][37] = 4;
        pixel_data[13][38] = 4;
        pixel_data[13][39] = 4;
        pixel_data[13][40] = 4;
        pixel_data[13][41] = 3;
        pixel_data[13][42] = 6;
        pixel_data[13][43] = 10;
        pixel_data[13][44] = 14;
        pixel_data[13][45] = 14;
        pixel_data[13][46] = 0;
        pixel_data[13][47] = 5;
        pixel_data[13][48] = 0;
        pixel_data[13][49] = 0; // y=13
        pixel_data[14][0] = 0;
        pixel_data[14][1] = 0;
        pixel_data[14][2] = 0;
        pixel_data[14][3] = 0;
        pixel_data[14][4] = 11;
        pixel_data[14][5] = 0;
        pixel_data[14][6] = 10;
        pixel_data[14][7] = 6;
        pixel_data[14][8] = 3;
        pixel_data[14][9] = 5;
        pixel_data[14][10] = 15;
        pixel_data[14][11] = 15;
        pixel_data[14][12] = 3;
        pixel_data[14][13] = 4;
        pixel_data[14][14] = 4;
        pixel_data[14][15] = 4;
        pixel_data[14][16] = 4;
        pixel_data[14][17] = 4;
        pixel_data[14][18] = 4;
        pixel_data[14][19] = 4;
        pixel_data[14][20] = 4;
        pixel_data[14][21] = 4;
        pixel_data[14][22] = 4;
        pixel_data[14][23] = 4;
        pixel_data[14][24] = 4;
        pixel_data[14][25] = 4;
        pixel_data[14][26] = 4;
        pixel_data[14][27] = 4;
        pixel_data[14][28] = 4;
        pixel_data[14][29] = 4;
        pixel_data[14][30] = 4;
        pixel_data[14][31] = 4;
        pixel_data[14][32] = 4;
        pixel_data[14][33] = 4;
        pixel_data[14][34] = 4;
        pixel_data[14][35] = 4;
        pixel_data[14][36] = 4;
        pixel_data[14][37] = 4;
        pixel_data[14][38] = 4;
        pixel_data[14][39] = 4;
        pixel_data[14][40] = 4;
        pixel_data[14][41] = 4;
        pixel_data[14][42] = 15;
        pixel_data[14][43] = 9;
        pixel_data[14][44] = 15;
        pixel_data[14][45] = 14;
        pixel_data[14][46] = 10;
        pixel_data[14][47] = 0;
        pixel_data[14][48] = 0;
        pixel_data[14][49] = 0; // y=14
        pixel_data[15][0] = 0;
        pixel_data[15][1] = 0;
        pixel_data[15][2] = 0;
        pixel_data[15][3] = 11;
        pixel_data[15][4] = 0;
        pixel_data[15][5] = 10;
        pixel_data[15][6] = 9;
        pixel_data[15][7] = 15;
        pixel_data[15][8] = 4;
        pixel_data[15][9] = 4;
        pixel_data[15][10] = 3;
        pixel_data[15][11] = 4;
        pixel_data[15][12] = 4;
        pixel_data[15][13] = 4;
        pixel_data[15][14] = 4;
        pixel_data[15][15] = 4;
        pixel_data[15][16] = 4;
        pixel_data[15][17] = 4;
        pixel_data[15][18] = 4;
        pixel_data[15][19] = 4;
        pixel_data[15][20] = 4;
        pixel_data[15][21] = 4;
        pixel_data[15][22] = 4;
        pixel_data[15][23] = 4;
        pixel_data[15][24] = 4;
        pixel_data[15][25] = 4;
        pixel_data[15][26] = 4;
        pixel_data[15][27] = 4;
        pixel_data[15][28] = 4;
        pixel_data[15][29] = 4;
        pixel_data[15][30] = 4;
        pixel_data[15][31] = 4;
        pixel_data[15][32] = 4;
        pixel_data[15][33] = 4;
        pixel_data[15][34] = 4;
        pixel_data[15][35] = 4;
        pixel_data[15][36] = 4;
        pixel_data[15][37] = 4;
        pixel_data[15][38] = 4;
        pixel_data[15][39] = 4;
        pixel_data[15][40] = 4;
        pixel_data[15][41] = 4;
        pixel_data[15][42] = 3;
        pixel_data[15][43] = 4;
        pixel_data[15][44] = 10;
        pixel_data[15][45] = 14;
        pixel_data[15][46] = 14;
        pixel_data[15][47] = 0;
        pixel_data[15][48] = 1;
        pixel_data[15][49] = 0; // y=15
        pixel_data[16][0] = 0;
        pixel_data[16][1] = 0;
        pixel_data[16][2] = 0;
        pixel_data[16][3] = 11;
        pixel_data[16][4] = 0;
        pixel_data[16][5] = 10;
        pixel_data[16][6] = 6;
        pixel_data[16][7] = 15;
        pixel_data[16][8] = 5;
        pixel_data[16][9] = 4;
        pixel_data[16][10] = 4;
        pixel_data[16][11] = 4;
        pixel_data[16][12] = 4;
        pixel_data[16][13] = 4;
        pixel_data[16][14] = 4;
        pixel_data[16][15] = 4;
        pixel_data[16][16] = 4;
        pixel_data[16][17] = 4;
        pixel_data[16][18] = 4;
        pixel_data[16][19] = 4;
        pixel_data[16][20] = 4;
        pixel_data[16][21] = 4;
        pixel_data[16][22] = 4;
        pixel_data[16][23] = 4;
        pixel_data[16][24] = 4;
        pixel_data[16][25] = 3;
        pixel_data[16][26] = 3;
        pixel_data[16][27] = 15;
        pixel_data[16][28] = 15;
        pixel_data[16][29] = 3;
        pixel_data[16][30] = 4;
        pixel_data[16][31] = 4;
        pixel_data[16][32] = 4;
        pixel_data[16][33] = 4;
        pixel_data[16][34] = 4;
        pixel_data[16][35] = 3;
        pixel_data[16][36] = 3;
        pixel_data[16][37] = 3;
        pixel_data[16][38] = 3;
        pixel_data[16][39] = 4;
        pixel_data[16][40] = 4;
        pixel_data[16][41] = 4;
        pixel_data[16][42] = 4;
        pixel_data[16][43] = 15;
        pixel_data[16][44] = 9;
        pixel_data[16][45] = 9;
        pixel_data[16][46] = 14;
        pixel_data[16][47] = 0;
        pixel_data[16][48] = 5;
        pixel_data[16][49] = 0; // y=16
        pixel_data[17][0] = 0;
        pixel_data[17][1] = 0;
        pixel_data[17][2] = 5;
        pixel_data[17][3] = 0;
        pixel_data[17][4] = 15;
        pixel_data[17][5] = 10;
        pixel_data[17][6] = 15;
        pixel_data[17][7] = 15;
        pixel_data[17][8] = 15;
        pixel_data[17][9] = 15;
        pixel_data[17][10] = 4;
        pixel_data[17][11] = 4;
        pixel_data[17][12] = 4;
        pixel_data[17][13] = 4;
        pixel_data[17][14] = 4;
        pixel_data[17][15] = 4;
        pixel_data[17][16] = 4;
        pixel_data[17][17] = 4;
        pixel_data[17][18] = 4;
        pixel_data[17][19] = 4;
        pixel_data[17][20] = 4;
        pixel_data[17][21] = 4;
        pixel_data[17][22] = 4;
        pixel_data[17][23] = 4;
        pixel_data[17][24] = 3;
        pixel_data[17][25] = 6;
        pixel_data[17][26] = 10;
        pixel_data[17][27] = 12;
        pixel_data[17][28] = 12;
        pixel_data[17][29] = 9;
        pixel_data[17][30] = 3;
        pixel_data[17][31] = 4;
        pixel_data[17][32] = 4;
        pixel_data[17][33] = 4;
        pixel_data[17][34] = 4;
        pixel_data[17][35] = 4;
        pixel_data[17][36] = 9;
        pixel_data[17][37] = 9;
        pixel_data[17][38] = 6;
        pixel_data[17][39] = 4;
        pixel_data[17][40] = 4;
        pixel_data[17][41] = 4;
        pixel_data[17][42] = 4;
        pixel_data[17][43] = 4;
        pixel_data[17][44] = 15;
        pixel_data[17][45] = 9;
        pixel_data[17][46] = 14;
        pixel_data[17][47] = 14;
        pixel_data[17][48] = 0;
        pixel_data[17][49] = 2; // y=17
        pixel_data[18][0] = 0;
        pixel_data[18][1] = 0;
        pixel_data[18][2] = 7;
        pixel_data[18][3] = 0;
        pixel_data[18][4] = 10;
        pixel_data[18][5] = 9;
        pixel_data[18][6] = 15;
        pixel_data[18][7] = 15;
        pixel_data[18][8] = 15;
        pixel_data[18][9] = 15;
        pixel_data[18][10] = 4;
        pixel_data[18][11] = 4;
        pixel_data[18][12] = 4;
        pixel_data[18][13] = 4;
        pixel_data[18][14] = 4;
        pixel_data[18][15] = 4;
        pixel_data[18][16] = 4;
        pixel_data[18][17] = 4;
        pixel_data[18][18] = 4;
        pixel_data[18][19] = 4;
        pixel_data[18][20] = 4;
        pixel_data[18][21] = 4;
        pixel_data[18][22] = 4;
        pixel_data[18][23] = 3;
        pixel_data[18][24] = 6;
        pixel_data[18][25] = 12;
        pixel_data[18][26] = 12;
        pixel_data[18][27] = 12;
        pixel_data[18][28] = 12;
        pixel_data[18][29] = 12;
        pixel_data[18][30] = 9;
        pixel_data[18][31] = 15;
        pixel_data[18][32] = 4;
        pixel_data[18][33] = 4;
        pixel_data[18][34] = 15;
        pixel_data[18][35] = 10;
        pixel_data[18][36] = 12;
        pixel_data[18][37] = 12;
        pixel_data[18][38] = 12;
        pixel_data[18][39] = 9;
        pixel_data[18][40] = 15;
        pixel_data[18][41] = 4;
        pixel_data[18][42] = 4;
        pixel_data[18][43] = 4;
        pixel_data[18][44] = 3;
        pixel_data[18][45] = 6;
        pixel_data[18][46] = 15;
        pixel_data[18][47] = 14;
        pixel_data[18][48] = 0;
        pixel_data[18][49] = 1; // y=18
        pixel_data[19][0] = 0;
        pixel_data[19][1] = 0;
        pixel_data[19][2] = 2;
        pixel_data[19][3] = 0;
        pixel_data[19][4] = 10;
        pixel_data[19][5] = 6;
        pixel_data[19][6] = 15;
        pixel_data[19][7] = 15;
        pixel_data[19][8] = 15;
        pixel_data[19][9] = 3;
        pixel_data[19][10] = 4;
        pixel_data[19][11] = 4;
        pixel_data[19][12] = 4;
        pixel_data[19][13] = 4;
        pixel_data[19][14] = 4;
        pixel_data[19][15] = 4;
        pixel_data[19][16] = 4;
        pixel_data[19][17] = 4;
        pixel_data[19][18] = 4;
        pixel_data[19][19] = 4;
        pixel_data[19][20] = 4;
        pixel_data[19][21] = 4;
        pixel_data[19][22] = 3;
        pixel_data[19][23] = 4;
        pixel_data[19][24] = 10;
        pixel_data[19][25] = 12;
        pixel_data[19][26] = 12;
        pixel_data[19][27] = 12;
        pixel_data[19][28] = 12;
        pixel_data[19][29] = 12;
        pixel_data[19][30] = 10;
        pixel_data[19][31] = 3;
        pixel_data[19][32] = 4;
        pixel_data[19][33] = 3;
        pixel_data[19][34] = 9;
        pixel_data[19][35] = 12;
        pixel_data[19][36] = 12;
        pixel_data[19][37] = 12;
        pixel_data[19][38] = 12;
        pixel_data[19][39] = 12;
        pixel_data[19][40] = 6;
        pixel_data[19][41] = 3;
        pixel_data[19][42] = 4;
        pixel_data[19][43] = 4;
        pixel_data[19][44] = 3;
        pixel_data[19][45] = 4;
        pixel_data[19][46] = 10;
        pixel_data[19][47] = 14;
        pixel_data[19][48] = 0;
        pixel_data[19][49] = 11; // y=19
        pixel_data[20][0] = 0;
        pixel_data[20][1] = 2;
        pixel_data[20][2] = 0;
        pixel_data[20][3] = 2;
        pixel_data[20][4] = 10;
        pixel_data[20][5] = 15;
        pixel_data[20][6] = 15;
        pixel_data[20][7] = 15;
        pixel_data[20][8] = 15;
        pixel_data[20][9] = 3;
        pixel_data[20][10] = 4;
        pixel_data[20][11] = 4;
        pixel_data[20][12] = 4;
        pixel_data[20][13] = 4;
        pixel_data[20][14] = 4;
        pixel_data[20][15] = 4;
        pixel_data[20][16] = 4;
        pixel_data[20][17] = 4;
        pixel_data[20][18] = 4;
        pixel_data[20][19] = 4;
        pixel_data[20][20] = 4;
        pixel_data[20][21] = 4;
        pixel_data[20][22] = 15;
        pixel_data[20][23] = 10;
        pixel_data[20][24] = 12;
        pixel_data[20][25] = 12;
        pixel_data[20][26] = 12;
        pixel_data[20][27] = 12;
        pixel_data[20][28] = 12;
        pixel_data[20][29] = 12;
        pixel_data[20][30] = 12;
        pixel_data[20][31] = 6;
        pixel_data[20][32] = 4;
        pixel_data[20][33] = 15;
        pixel_data[20][34] = 10;
        pixel_data[20][35] = 12;
        pixel_data[20][36] = 12;
        pixel_data[20][37] = 12;
        pixel_data[20][38] = 12;
        pixel_data[20][39] = 2;
        pixel_data[20][40] = 10;
        pixel_data[20][41] = 15;
        pixel_data[20][42] = 4;
        pixel_data[20][43] = 4;
        pixel_data[20][44] = 4;
        pixel_data[20][45] = 15;
        pixel_data[20][46] = 9;
        pixel_data[20][47] = 10;
        pixel_data[20][48] = 0;
        pixel_data[20][49] = 2; // y=20
        pixel_data[21][0] = 0;
        pixel_data[21][1] = 10;
        pixel_data[21][2] = 0;
        pixel_data[21][3] = 12;
        pixel_data[21][4] = 9;
        pixel_data[21][5] = 15;
        pixel_data[21][6] = 15;
        pixel_data[21][7] = 15;
        pixel_data[21][8] = 15;
        pixel_data[21][9] = 4;
        pixel_data[21][10] = 4;
        pixel_data[21][11] = 4;
        pixel_data[21][12] = 4;
        pixel_data[21][13] = 4;
        pixel_data[21][14] = 4;
        pixel_data[21][15] = 4;
        pixel_data[21][16] = 4;
        pixel_data[21][17] = 4;
        pixel_data[21][18] = 4;
        pixel_data[21][19] = 4;
        pixel_data[21][20] = 4;
        pixel_data[21][21] = 4;
        pixel_data[21][22] = 3;
        pixel_data[21][23] = 12;
        pixel_data[21][24] = 12;
        pixel_data[21][25] = 12;
        pixel_data[21][26] = 12;
        pixel_data[21][27] = 12;
        pixel_data[21][28] = 12;
        pixel_data[21][29] = 12;
        pixel_data[21][30] = 12;
        pixel_data[21][31] = 9;
        pixel_data[21][32] = 3;
        pixel_data[21][33] = 15;
        pixel_data[21][34] = 9;
        pixel_data[21][35] = 12;
        pixel_data[21][36] = 12;
        pixel_data[21][37] = 12;
        pixel_data[21][38] = 12;
        pixel_data[21][39] = 12;
        pixel_data[21][40] = 12;
        pixel_data[21][41] = 4;
        pixel_data[21][42] = 4;
        pixel_data[21][43] = 4;
        pixel_data[21][44] = 4;
        pixel_data[21][45] = 15;
        pixel_data[21][46] = 6;
        pixel_data[21][47] = 10;
        pixel_data[21][48] = 5;
        pixel_data[21][49] = 0; // y=21
        pixel_data[22][0] = 0;
        pixel_data[22][1] = 11;
        pixel_data[22][2] = 0;
        pixel_data[22][3] = 11;
        pixel_data[22][4] = 6;
        pixel_data[22][5] = 15;
        pixel_data[22][6] = 15;
        pixel_data[22][7] = 15;
        pixel_data[22][8] = 15;
        pixel_data[22][9] = 4;
        pixel_data[22][10] = 4;
        pixel_data[22][11] = 4;
        pixel_data[22][12] = 4;
        pixel_data[22][13] = 4;
        pixel_data[22][14] = 4;
        pixel_data[22][15] = 4;
        pixel_data[22][16] = 4;
        pixel_data[22][17] = 4;
        pixel_data[22][18] = 4;
        pixel_data[22][19] = 4;
        pixel_data[22][20] = 4;
        pixel_data[22][21] = 4;
        pixel_data[22][22] = 3;
        pixel_data[22][23] = 10;
        pixel_data[22][24] = 12;
        pixel_data[22][25] = 12;
        pixel_data[22][26] = 12;
        pixel_data[22][27] = 12;
        pixel_data[22][28] = 12;
        pixel_data[22][29] = 12;
        pixel_data[22][30] = 12;
        pixel_data[22][31] = 9;
        pixel_data[22][32] = 3;
        pixel_data[22][33] = 3;
        pixel_data[22][34] = 6;
        pixel_data[22][35] = 12;
        pixel_data[22][36] = 12;
        pixel_data[22][37] = 12;
        pixel_data[22][38] = 12;
        pixel_data[22][39] = 12;
        pixel_data[22][40] = 12;
        pixel_data[22][41] = 6;
        pixel_data[22][42] = 3;
        pixel_data[22][43] = 4;
        pixel_data[22][44] = 4;
        pixel_data[22][45] = 4;
        pixel_data[22][46] = 3;
        pixel_data[22][47] = 10;
        pixel_data[22][48] = 10;
        pixel_data[22][49] = 0; // y=22
        pixel_data[23][0] = 2;
        pixel_data[23][1] = 0;
        pixel_data[23][2] = 2;
        pixel_data[23][3] = 11;
        pixel_data[23][4] = 3;
        pixel_data[23][5] = 15;
        pixel_data[23][6] = 15;
        pixel_data[23][7] = 15;
        pixel_data[23][8] = 15;
        pixel_data[23][9] = 4;
        pixel_data[23][10] = 4;
        pixel_data[23][11] = 4;
        pixel_data[23][12] = 4;
        pixel_data[23][13] = 4;
        pixel_data[23][14] = 4;
        pixel_data[23][15] = 4;
        pixel_data[23][16] = 4;
        pixel_data[23][17] = 4;
        pixel_data[23][18] = 4;
        pixel_data[23][19] = 4;
        pixel_data[23][20] = 4;
        pixel_data[23][21] = 4;
        pixel_data[23][22] = 15;
        pixel_data[23][23] = 10;
        pixel_data[23][24] = 12;
        pixel_data[23][25] = 12;
        pixel_data[23][26] = 12;
        pixel_data[23][27] = 12;
        pixel_data[23][28] = 12;
        pixel_data[23][29] = 12;
        pixel_data[23][30] = 12;
        pixel_data[23][31] = 6;
        pixel_data[23][32] = 3;
        pixel_data[23][33] = 4;
        pixel_data[23][34] = 3;
        pixel_data[23][35] = 12;
        pixel_data[23][36] = 12;
        pixel_data[23][37] = 12;
        pixel_data[23][38] = 12;
        pixel_data[23][39] = 12;
        pixel_data[23][40] = 12;
        pixel_data[23][41] = 4;
        pixel_data[23][42] = 3;
        pixel_data[23][43] = 4;
        pixel_data[23][44] = 4;
        pixel_data[23][45] = 4;
        pixel_data[23][46] = 3;
        pixel_data[23][47] = 9;
        pixel_data[23][48] = 12;
        pixel_data[23][49] = 0; // y=23
        pixel_data[24][0] = 13;
        pixel_data[24][1] = 0;
        pixel_data[24][2] = 2;
        pixel_data[24][3] = 11;
        pixel_data[24][4] = 15;
        pixel_data[24][5] = 15;
        pixel_data[24][6] = 15;
        pixel_data[24][7] = 15;
        pixel_data[24][8] = 4;
        pixel_data[24][9] = 4;
        pixel_data[24][10] = 4;
        pixel_data[24][11] = 4;
        pixel_data[24][12] = 4;
        pixel_data[24][13] = 4;
        pixel_data[24][14] = 4;
        pixel_data[24][15] = 4;
        pixel_data[24][16] = 4;
        pixel_data[24][17] = 4;
        pixel_data[24][18] = 4;
        pixel_data[24][19] = 4;
        pixel_data[24][20] = 4;
        pixel_data[24][21] = 4;
        pixel_data[24][22] = 3;
        pixel_data[24][23] = 6;
        pixel_data[24][24] = 12;
        pixel_data[24][25] = 12;
        pixel_data[24][26] = 12;
        pixel_data[24][27] = 12;
        pixel_data[24][28] = 12;
        pixel_data[24][29] = 12;
        pixel_data[24][30] = 10;
        pixel_data[24][31] = 3;
        pixel_data[24][32] = 4;
        pixel_data[24][33] = 4;
        pixel_data[24][34] = 15;
        pixel_data[24][35] = 9;
        pixel_data[24][36] = 12;
        pixel_data[24][37] = 12;
        pixel_data[24][38] = 12;
        pixel_data[24][39] = 2;
        pixel_data[24][40] = 10;
        pixel_data[24][41] = 15;
        pixel_data[24][42] = 4;
        pixel_data[24][43] = 4;
        pixel_data[24][44] = 4;
        pixel_data[24][45] = 4;
        pixel_data[24][46] = 3;
        pixel_data[24][47] = 3;
        pixel_data[24][48] = 13;
        pixel_data[24][49] = 0; // y=24
        pixel_data[25][0] = 11;
        pixel_data[25][1] = 0;
        pixel_data[25][2] = 1;
        pixel_data[25][3] = 5;
        pixel_data[25][4] = 3;
        pixel_data[25][5] = 3;
        pixel_data[25][6] = 15;
        pixel_data[25][7] = 4;
        pixel_data[25][8] = 4;
        pixel_data[25][9] = 4;
        pixel_data[25][10] = 4;
        pixel_data[25][11] = 4;
        pixel_data[25][12] = 4;
        pixel_data[25][13] = 4;
        pixel_data[25][14] = 4;
        pixel_data[25][15] = 4;
        pixel_data[25][16] = 4;
        pixel_data[25][17] = 4;
        pixel_data[25][18] = 4;
        pixel_data[25][19] = 4;
        pixel_data[25][20] = 4;
        pixel_data[25][21] = 4;
        pixel_data[25][22] = 4;
        pixel_data[25][23] = 3;
        pixel_data[25][24] = 9;
        pixel_data[25][25] = 10;
        pixel_data[25][26] = 12;
        pixel_data[25][27] = 12;
        pixel_data[25][28] = 12;
        pixel_data[25][29] = 12;
        pixel_data[25][30] = 9;
        pixel_data[25][31] = 3;
        pixel_data[25][32] = 4;
        pixel_data[25][33] = 4;
        pixel_data[25][34] = 4;
        pixel_data[25][35] = 4;
        pixel_data[25][36] = 9;
        pixel_data[25][37] = 9;
        pixel_data[25][38] = 10;
        pixel_data[25][39] = 9;
        pixel_data[25][40] = 6;
        pixel_data[25][41] = 3;
        pixel_data[25][42] = 4;
        pixel_data[25][43] = 4;
        pixel_data[25][44] = 4;
        pixel_data[25][45] = 4;
        pixel_data[25][46] = 4;
        pixel_data[25][47] = 15;
        pixel_data[25][48] = 11;
        pixel_data[25][49] = 2; // y=25
        pixel_data[26][0] = 6;
        pixel_data[26][1] = 0;
        pixel_data[26][2] = 13;
        pixel_data[26][3] = 15;
        pixel_data[26][4] = 4;
        pixel_data[26][5] = 4;
        pixel_data[26][6] = 4;
        pixel_data[26][7] = 4;
        pixel_data[26][8] = 4;
        pixel_data[26][9] = 4;
        pixel_data[26][10] = 4;
        pixel_data[26][11] = 4;
        pixel_data[26][12] = 4;
        pixel_data[26][13] = 4;
        pixel_data[26][14] = 4;
        pixel_data[26][15] = 4;
        pixel_data[26][16] = 4;
        pixel_data[26][17] = 4;
        pixel_data[26][18] = 4;
        pixel_data[26][19] = 4;
        pixel_data[26][20] = 4;
        pixel_data[26][21] = 4;
        pixel_data[26][22] = 4;
        pixel_data[26][23] = 4;
        pixel_data[26][24] = 3;
        pixel_data[26][25] = 4;
        pixel_data[26][26] = 6;
        pixel_data[26][27] = 10;
        pixel_data[26][28] = 10;
        pixel_data[26][29] = 6;
        pixel_data[26][30] = 3;
        pixel_data[26][31] = 4;
        pixel_data[26][32] = 4;
        pixel_data[26][33] = 4;
        pixel_data[26][34] = 4;
        pixel_data[26][35] = 4;
        pixel_data[26][36] = 15;
        pixel_data[26][37] = 15;
        pixel_data[26][38] = 3;
        pixel_data[26][39] = 3;
        pixel_data[26][40] = 3;
        pixel_data[26][41] = 4;
        pixel_data[26][42] = 4;
        pixel_data[26][43] = 4;
        pixel_data[26][44] = 4;
        pixel_data[26][45] = 4;
        pixel_data[26][46] = 4;
        pixel_data[26][47] = 15;
        pixel_data[26][48] = 11;
        pixel_data[26][49] = 2; // y=26
        pixel_data[27][0] = 0;
        pixel_data[27][1] = 2;
        pixel_data[27][2] = 11;
        pixel_data[27][3] = 15;
        pixel_data[27][4] = 4;
        pixel_data[27][5] = 4;
        pixel_data[27][6] = 4;
        pixel_data[27][7] = 4;
        pixel_data[27][8] = 4;
        pixel_data[27][9] = 4;
        pixel_data[27][10] = 4;
        pixel_data[27][11] = 4;
        pixel_data[27][12] = 4;
        pixel_data[27][13] = 4;
        pixel_data[27][14] = 4;
        pixel_data[27][15] = 4;
        pixel_data[27][16] = 4;
        pixel_data[27][17] = 4;
        pixel_data[27][18] = 4;
        pixel_data[27][19] = 4;
        pixel_data[27][20] = 4;
        pixel_data[27][21] = 4;
        pixel_data[27][22] = 4;
        pixel_data[27][23] = 4;
        pixel_data[27][24] = 4;
        pixel_data[27][25] = 4;
        pixel_data[27][26] = 3;
        pixel_data[27][27] = 4;
        pixel_data[27][28] = 4;
        pixel_data[27][29] = 3;
        pixel_data[27][30] = 4;
        pixel_data[27][31] = 4;
        pixel_data[27][32] = 4;
        pixel_data[27][33] = 3;
        pixel_data[27][34] = 4;
        pixel_data[27][35] = 4;
        pixel_data[27][36] = 4;
        pixel_data[27][37] = 4;
        pixel_data[27][38] = 4;
        pixel_data[27][39] = 4;
        pixel_data[27][40] = 4;
        pixel_data[27][41] = 4;
        pixel_data[27][42] = 4;
        pixel_data[27][43] = 4;
        pixel_data[27][44] = 4;
        pixel_data[27][45] = 4;
        pixel_data[27][46] = 4;
        pixel_data[27][47] = 3;
        pixel_data[27][48] = 11;
        pixel_data[27][49] = 1; // y=27
        pixel_data[28][0] = 0;
        pixel_data[28][1] = 2;
        pixel_data[28][2] = 11;
        pixel_data[28][3] = 15;
        pixel_data[28][4] = 4;
        pixel_data[28][5] = 4;
        pixel_data[28][6] = 4;
        pixel_data[28][7] = 4;
        pixel_data[28][8] = 4;
        pixel_data[28][9] = 4;
        pixel_data[28][10] = 4;
        pixel_data[28][11] = 4;
        pixel_data[28][12] = 4;
        pixel_data[28][13] = 4;
        pixel_data[28][14] = 4;
        pixel_data[28][15] = 4;
        pixel_data[28][16] = 4;
        pixel_data[28][17] = 4;
        pixel_data[28][18] = 4;
        pixel_data[28][19] = 4;
        pixel_data[28][20] = 4;
        pixel_data[28][21] = 4;
        pixel_data[28][22] = 4;
        pixel_data[28][23] = 4;
        pixel_data[28][24] = 4;
        pixel_data[28][25] = 4;
        pixel_data[28][26] = 4;
        pixel_data[28][27] = 3;
        pixel_data[28][28] = 3;
        pixel_data[28][29] = 4;
        pixel_data[28][30] = 4;
        pixel_data[28][31] = 3;
        pixel_data[28][32] = 4;
        pixel_data[28][33] = 9;
        pixel_data[28][34] = 15;
        pixel_data[28][35] = 4;
        pixel_data[28][36] = 4;
        pixel_data[28][37] = 4;
        pixel_data[28][38] = 4;
        pixel_data[28][39] = 4;
        pixel_data[28][40] = 4;
        pixel_data[28][41] = 4;
        pixel_data[28][42] = 4;
        pixel_data[28][43] = 4;
        pixel_data[28][44] = 4;
        pixel_data[28][45] = 4;
        pixel_data[28][46] = 4;
        pixel_data[28][47] = 5;
        pixel_data[28][48] = 8;
        pixel_data[28][49] = 1; // y=28
        pixel_data[29][0] = 0;
        pixel_data[29][1] = 1;
        pixel_data[29][2] = 11;
        pixel_data[29][3] = 15;
        pixel_data[29][4] = 4;
        pixel_data[29][5] = 4;
        pixel_data[29][6] = 4;
        pixel_data[29][7] = 4;
        pixel_data[29][8] = 4;
        pixel_data[29][9] = 4;
        pixel_data[29][10] = 4;
        pixel_data[29][11] = 4;
        pixel_data[29][12] = 4;
        pixel_data[29][13] = 4;
        pixel_data[29][14] = 4;
        pixel_data[29][15] = 4;
        pixel_data[29][16] = 4;
        pixel_data[29][17] = 4;
        pixel_data[29][18] = 4;
        pixel_data[29][19] = 4;
        pixel_data[29][20] = 4;
        pixel_data[29][21] = 4;
        pixel_data[29][22] = 4;
        pixel_data[29][23] = 4;
        pixel_data[29][24] = 4;
        pixel_data[29][25] = 4;
        pixel_data[29][26] = 4;
        pixel_data[29][27] = 4;
        pixel_data[29][28] = 4;
        pixel_data[29][29] = 4;
        pixel_data[29][30] = 3;
        pixel_data[29][31] = 6;
        pixel_data[29][32] = 10;
        pixel_data[29][33] = 12;
        pixel_data[29][34] = 10;
        pixel_data[29][35] = 4;
        pixel_data[29][36] = 3;
        pixel_data[29][37] = 4;
        pixel_data[29][38] = 4;
        pixel_data[29][39] = 4;
        pixel_data[29][40] = 4;
        pixel_data[29][41] = 4;
        pixel_data[29][42] = 4;
        pixel_data[29][43] = 4;
        pixel_data[29][44] = 4;
        pixel_data[29][45] = 4;
        pixel_data[29][46] = 4;
        pixel_data[29][47] = 5;
        pixel_data[29][48] = 8;
        pixel_data[29][49] = 13; // y=29
        pixel_data[30][0] = 0;
        pixel_data[30][1] = 1;
        pixel_data[30][2] = 8;
        pixel_data[30][3] = 15;
        pixel_data[30][4] = 6;
        pixel_data[30][5] = 4;
        pixel_data[30][6] = 4;
        pixel_data[30][7] = 4;
        pixel_data[30][8] = 4;
        pixel_data[30][9] = 4;
        pixel_data[30][10] = 4;
        pixel_data[30][11] = 4;
        pixel_data[30][12] = 4;
        pixel_data[30][13] = 4;
        pixel_data[30][14] = 4;
        pixel_data[30][15] = 4;
        pixel_data[30][16] = 4;
        pixel_data[30][17] = 4;
        pixel_data[30][18] = 4;
        pixel_data[30][19] = 4;
        pixel_data[30][20] = 4;
        pixel_data[30][21] = 4;
        pixel_data[30][22] = 4;
        pixel_data[30][23] = 4;
        pixel_data[30][24] = 4;
        pixel_data[30][25] = 4;
        pixel_data[30][26] = 4;
        pixel_data[30][27] = 4;
        pixel_data[30][28] = 4;
        pixel_data[30][29] = 3;
        pixel_data[30][30] = 6;
        pixel_data[30][31] = 12;
        pixel_data[30][32] = 12;
        pixel_data[30][33] = 12;
        pixel_data[30][34] = 12;
        pixel_data[30][35] = 10;
        pixel_data[30][36] = 15;
        pixel_data[30][37] = 4;
        pixel_data[30][38] = 4;
        pixel_data[30][39] = 4;
        pixel_data[30][40] = 4;
        pixel_data[30][41] = 4;
        pixel_data[30][42] = 4;
        pixel_data[30][43] = 4;
        pixel_data[30][44] = 4;
        pixel_data[30][45] = 4;
        pixel_data[30][46] = 4;
        pixel_data[30][47] = 5;
        pixel_data[30][48] = 8;
        pixel_data[30][49] = 11; // y=30
        pixel_data[31][0] = 0;
        pixel_data[31][1] = 1;
        pixel_data[31][2] = 8;
        pixel_data[31][3] = 8;
        pixel_data[31][4] = 6;
        pixel_data[31][5] = 4;
        pixel_data[31][6] = 4;
        pixel_data[31][7] = 4;
        pixel_data[31][8] = 4;
        pixel_data[31][9] = 4;
        pixel_data[31][10] = 4;
        pixel_data[31][11] = 4;
        pixel_data[31][12] = 4;
        pixel_data[31][13] = 4;
        pixel_data[31][14] = 4;
        pixel_data[31][15] = 4;
        pixel_data[31][16] = 4;
        pixel_data[31][17] = 4;
        pixel_data[31][18] = 4;
        pixel_data[31][19] = 4;
        pixel_data[31][20] = 4;
        pixel_data[31][21] = 4;
        pixel_data[31][22] = 4;
        pixel_data[31][23] = 4;
        pixel_data[31][24] = 4;
        pixel_data[31][25] = 4;
        pixel_data[31][26] = 4;
        pixel_data[31][27] = 4;
        pixel_data[31][28] = 4;
        pixel_data[31][29] = 15;
        pixel_data[31][30] = 9;
        pixel_data[31][31] = 12;
        pixel_data[31][32] = 12;
        pixel_data[31][33] = 12;
        pixel_data[31][34] = 12;
        pixel_data[31][35] = 12;
        pixel_data[31][36] = 6;
        pixel_data[31][37] = 3;
        pixel_data[31][38] = 4;
        pixel_data[31][39] = 4;
        pixel_data[31][40] = 4;
        pixel_data[31][41] = 4;
        pixel_data[31][42] = 4;
        pixel_data[31][43] = 4;
        pixel_data[31][44] = 4;
        pixel_data[31][45] = 4;
        pixel_data[31][46] = 3;
        pixel_data[31][47] = 8;
        pixel_data[31][48] = 8;
        pixel_data[31][49] = 11; // y=31
        pixel_data[32][0] = 0;
        pixel_data[32][1] = 1;
        pixel_data[32][2] = 8;
        pixel_data[32][3] = 8;
        pixel_data[32][4] = 5;
        pixel_data[32][5] = 4;
        pixel_data[32][6] = 4;
        pixel_data[32][7] = 4;
        pixel_data[32][8] = 4;
        pixel_data[32][9] = 4;
        pixel_data[32][10] = 4;
        pixel_data[32][11] = 4;
        pixel_data[32][12] = 4;
        pixel_data[32][13] = 4;
        pixel_data[32][14] = 4;
        pixel_data[32][15] = 4;
        pixel_data[32][16] = 4;
        pixel_data[32][17] = 4;
        pixel_data[32][18] = 4;
        pixel_data[32][19] = 4;
        pixel_data[32][20] = 4;
        pixel_data[32][21] = 4;
        pixel_data[32][22] = 4;
        pixel_data[32][23] = 4;
        pixel_data[32][24] = 4;
        pixel_data[32][25] = 4;
        pixel_data[32][26] = 4;
        pixel_data[32][27] = 4;
        pixel_data[32][28] = 4;
        pixel_data[32][29] = 15;
        pixel_data[32][30] = 10;
        pixel_data[32][31] = 12;
        pixel_data[32][32] = 12;
        pixel_data[32][33] = 12;
        pixel_data[32][34] = 12;
        pixel_data[32][35] = 12;
        pixel_data[32][36] = 9;
        pixel_data[32][37] = 15;
        pixel_data[32][38] = 4;
        pixel_data[32][39] = 4;
        pixel_data[32][40] = 4;
        pixel_data[32][41] = 4;
        pixel_data[32][42] = 4;
        pixel_data[32][43] = 4;
        pixel_data[32][44] = 4;
        pixel_data[32][45] = 4;
        pixel_data[32][46] = 6;
        pixel_data[32][47] = 8;
        pixel_data[32][48] = 8;
        pixel_data[32][49] = 8; // y=32
        pixel_data[33][0] = 0;
        pixel_data[33][1] = 1;
        pixel_data[33][2] = 8;
        pixel_data[33][3] = 8;
        pixel_data[33][4] = 15;
        pixel_data[33][5] = 4;
        pixel_data[33][6] = 4;
        pixel_data[33][7] = 4;
        pixel_data[33][8] = 4;
        pixel_data[33][9] = 4;
        pixel_data[33][10] = 4;
        pixel_data[33][11] = 4;
        pixel_data[33][12] = 4;
        pixel_data[33][13] = 4;
        pixel_data[33][14] = 4;
        pixel_data[33][15] = 4;
        pixel_data[33][16] = 4;
        pixel_data[33][17] = 4;
        pixel_data[33][18] = 4;
        pixel_data[33][19] = 4;
        pixel_data[33][20] = 4;
        pixel_data[33][21] = 4;
        pixel_data[33][22] = 4;
        pixel_data[33][23] = 4;
        pixel_data[33][24] = 4;
        pixel_data[33][25] = 4;
        pixel_data[33][26] = 4;
        pixel_data[33][27] = 4;
        pixel_data[33][28] = 4;
        pixel_data[33][29] = 15;
        pixel_data[33][30] = 10;
        pixel_data[33][31] = 12;
        pixel_data[33][32] = 12;
        pixel_data[33][33] = 12;
        pixel_data[33][34] = 12;
        pixel_data[33][35] = 12;
        pixel_data[33][36] = 10;
        pixel_data[33][37] = 15;
        pixel_data[33][38] = 4;
        pixel_data[33][39] = 4;
        pixel_data[33][40] = 4;
        pixel_data[33][41] = 4;
        pixel_data[33][42] = 4;
        pixel_data[33][43] = 4;
        pixel_data[33][44] = 4;
        pixel_data[33][45] = 4;
        pixel_data[33][46] = 5;
        pixel_data[33][47] = 8;
        pixel_data[33][48] = 8;
        pixel_data[33][49] = 8; // y=33
        pixel_data[34][0] = 0;
        pixel_data[34][1] = 1;
        pixel_data[34][2] = 8;
        pixel_data[34][3] = 8;
        pixel_data[34][4] = 8;
        pixel_data[34][5] = 3;
        pixel_data[34][6] = 4;
        pixel_data[34][7] = 4;
        pixel_data[34][8] = 4;
        pixel_data[34][9] = 4;
        pixel_data[34][10] = 4;
        pixel_data[34][11] = 4;
        pixel_data[34][12] = 4;
        pixel_data[34][13] = 4;
        pixel_data[34][14] = 4;
        pixel_data[34][15] = 4;
        pixel_data[34][16] = 4;
        pixel_data[34][17] = 4;
        pixel_data[34][18] = 4;
        pixel_data[34][19] = 4;
        pixel_data[34][20] = 4;
        pixel_data[34][21] = 4;
        pixel_data[34][22] = 4;
        pixel_data[34][23] = 4;
        pixel_data[34][24] = 4;
        pixel_data[34][25] = 4;
        pixel_data[34][26] = 4;
        pixel_data[34][27] = 4;
        pixel_data[34][28] = 4;
        pixel_data[34][29] = 15;
        pixel_data[34][30] = 10;
        pixel_data[34][31] = 12;
        pixel_data[34][32] = 12;
        pixel_data[34][33] = 12;
        pixel_data[34][34] = 12;
        pixel_data[34][35] = 12;
        pixel_data[34][36] = 9;
        pixel_data[34][37] = 15;
        pixel_data[34][38] = 4;
        pixel_data[34][39] = 4;
        pixel_data[34][40] = 4;
        pixel_data[34][41] = 4;
        pixel_data[34][42] = 4;
        pixel_data[34][43] = 4;
        pixel_data[34][44] = 4;
        pixel_data[34][45] = 4;
        pixel_data[34][46] = 8;
        pixel_data[34][47] = 8;
        pixel_data[34][48] = 8;
        pixel_data[34][49] = 8; // y=34
        pixel_data[35][0] = 0;
        pixel_data[35][1] = 1;
        pixel_data[35][2] = 8;
        pixel_data[35][3] = 8;
        pixel_data[35][4] = 8;
        pixel_data[35][5] = 5;
        pixel_data[35][6] = 4;
        pixel_data[35][7] = 4;
        pixel_data[35][8] = 4;
        pixel_data[35][9] = 4;
        pixel_data[35][10] = 4;
        pixel_data[35][11] = 4;
        pixel_data[35][12] = 4;
        pixel_data[35][13] = 4;
        pixel_data[35][14] = 4;
        pixel_data[35][15] = 4;
        pixel_data[35][16] = 4;
        pixel_data[35][17] = 4;
        pixel_data[35][18] = 4;
        pixel_data[35][19] = 4;
        pixel_data[35][20] = 4;
        pixel_data[35][21] = 4;
        pixel_data[35][22] = 4;
        pixel_data[35][23] = 4;
        pixel_data[35][24] = 4;
        pixel_data[35][25] = 4;
        pixel_data[35][26] = 4;
        pixel_data[35][27] = 4;
        pixel_data[35][28] = 4;
        pixel_data[35][29] = 15;
        pixel_data[35][30] = 10;
        pixel_data[35][31] = 12;
        pixel_data[35][32] = 12;
        pixel_data[35][33] = 12;
        pixel_data[35][34] = 12;
        pixel_data[35][35] = 12;
        pixel_data[35][36] = 9;
        pixel_data[35][37] = 15;
        pixel_data[35][38] = 4;
        pixel_data[35][39] = 4;
        pixel_data[35][40] = 4;
        pixel_data[35][41] = 4;
        pixel_data[35][42] = 4;
        pixel_data[35][43] = 4;
        pixel_data[35][44] = 4;
        pixel_data[35][45] = 5;
        pixel_data[35][46] = 8;
        pixel_data[35][47] = 8;
        pixel_data[35][48] = 8;
        pixel_data[35][49] = 8; // y=35
        pixel_data[36][0] = 0;
        pixel_data[36][1] = 13;
        pixel_data[36][2] = 8;
        pixel_data[36][3] = 8;
        pixel_data[36][4] = 8;
        pixel_data[36][5] = 8;
        pixel_data[36][6] = 4;
        pixel_data[36][7] = 4;
        pixel_data[36][8] = 4;
        pixel_data[36][9] = 4;
        pixel_data[36][10] = 4;
        pixel_data[36][11] = 4;
        pixel_data[36][12] = 4;
        pixel_data[36][13] = 4;
        pixel_data[36][14] = 4;
        pixel_data[36][15] = 4;
        pixel_data[36][16] = 4;
        pixel_data[36][17] = 4;
        pixel_data[36][18] = 4;
        pixel_data[36][19] = 4;
        pixel_data[36][20] = 4;
        pixel_data[36][21] = 4;
        pixel_data[36][22] = 4;
        pixel_data[36][23] = 4;
        pixel_data[36][24] = 4;
        pixel_data[36][25] = 4;
        pixel_data[36][26] = 4;
        pixel_data[36][27] = 4;
        pixel_data[36][28] = 4;
        pixel_data[36][29] = 3;
        pixel_data[36][30] = 6;
        pixel_data[36][31] = 12;
        pixel_data[36][32] = 12;
        pixel_data[36][33] = 12;
        pixel_data[36][34] = 12;
        pixel_data[36][35] = 10;
        pixel_data[36][36] = 3;
        pixel_data[36][37] = 4;
        pixel_data[36][38] = 4;
        pixel_data[36][39] = 4;
        pixel_data[36][40] = 4;
        pixel_data[36][41] = 4;
        pixel_data[36][42] = 4;
        pixel_data[36][43] = 4;
        pixel_data[36][44] = 4;
        pixel_data[36][45] = 8;
        pixel_data[36][46] = 8;
        pixel_data[36][47] = 8;
        pixel_data[36][48] = 8;
        pixel_data[36][49] = 8; // y=36
        pixel_data[37][0] = 0;
        pixel_data[37][1] = 13;
        pixel_data[37][2] = 8;
        pixel_data[37][3] = 8;
        pixel_data[37][4] = 8;
        pixel_data[37][5] = 8;
        pixel_data[37][6] = 5;
        pixel_data[37][7] = 4;
        pixel_data[37][8] = 4;
        pixel_data[37][9] = 4;
        pixel_data[37][10] = 4;
        pixel_data[37][11] = 4;
        pixel_data[37][12] = 4;
        pixel_data[37][13] = 4;
        pixel_data[37][14] = 4;
        pixel_data[37][15] = 4;
        pixel_data[37][16] = 4;
        pixel_data[37][17] = 4;
        pixel_data[37][18] = 4;
        pixel_data[37][19] = 4;
        pixel_data[37][20] = 4;
        pixel_data[37][21] = 4;
        pixel_data[37][22] = 4;
        pixel_data[37][23] = 4;
        pixel_data[37][24] = 4;
        pixel_data[37][25] = 4;
        pixel_data[37][26] = 4;
        pixel_data[37][27] = 4;
        pixel_data[37][28] = 4;
        pixel_data[37][29] = 4;
        pixel_data[37][30] = 3;
        pixel_data[37][31] = 9;
        pixel_data[37][32] = 12;
        pixel_data[37][33] = 12;
        pixel_data[37][34] = 12;
        pixel_data[37][35] = 9;
        pixel_data[37][36] = 15;
        pixel_data[37][37] = 4;
        pixel_data[37][38] = 4;
        pixel_data[37][39] = 4;
        pixel_data[37][40] = 4;
        pixel_data[37][41] = 4;
        pixel_data[37][42] = 4;
        pixel_data[37][43] = 4;
        pixel_data[37][44] = 5;
        pixel_data[37][45] = 8;
        pixel_data[37][46] = 8;
        pixel_data[37][47] = 8;
        pixel_data[37][48] = 8;
        pixel_data[37][49] = 8; // y=37
        pixel_data[38][0] = 0;
        pixel_data[38][1] = 13;
        pixel_data[38][2] = 8;
        pixel_data[38][3] = 8;
        pixel_data[38][4] = 8;
        pixel_data[38][5] = 8;
        pixel_data[38][6] = 8;
        pixel_data[38][7] = 6;
        pixel_data[38][8] = 4;
        pixel_data[38][9] = 4;
        pixel_data[38][10] = 4;
        pixel_data[38][11] = 4;
        pixel_data[38][12] = 4;
        pixel_data[38][13] = 4;
        pixel_data[38][14] = 4;
        pixel_data[38][15] = 4;
        pixel_data[38][16] = 4;
        pixel_data[38][17] = 4;
        pixel_data[38][18] = 4;
        pixel_data[38][19] = 4;
        pixel_data[38][20] = 4;
        pixel_data[38][21] = 4;
        pixel_data[38][22] = 4;
        pixel_data[38][23] = 4;
        pixel_data[38][24] = 4;
        pixel_data[38][25] = 4;
        pixel_data[38][26] = 4;
        pixel_data[38][27] = 4;
        pixel_data[38][28] = 4;
        pixel_data[38][29] = 4;
        pixel_data[38][30] = 4;
        pixel_data[38][31] = 3;
        pixel_data[38][32] = 6;
        pixel_data[38][33] = 6;
        pixel_data[38][34] = 6;
        pixel_data[38][35] = 3;
        pixel_data[38][36] = 4;
        pixel_data[38][37] = 4;
        pixel_data[38][38] = 4;
        pixel_data[38][39] = 4;
        pixel_data[38][40] = 4;
        pixel_data[38][41] = 4;
        pixel_data[38][42] = 4;
        pixel_data[38][43] = 4;
        pixel_data[38][44] = 8;
        pixel_data[38][45] = 8;
        pixel_data[38][46] = 8;
        pixel_data[38][47] = 8;
        pixel_data[38][48] = 8;
        pixel_data[38][49] = 8; // y=38
        pixel_data[39][0] = 0;
        pixel_data[39][1] = 13;
        pixel_data[39][2] = 8;
        pixel_data[39][3] = 8;
        pixel_data[39][4] = 8;
        pixel_data[39][5] = 8;
        pixel_data[39][6] = 8;
        pixel_data[39][7] = 15;
        pixel_data[39][8] = 4;
        pixel_data[39][9] = 4;
        pixel_data[39][10] = 4;
        pixel_data[39][11] = 4;
        pixel_data[39][12] = 4;
        pixel_data[39][13] = 4;
        pixel_data[39][14] = 4;
        pixel_data[39][15] = 4;
        pixel_data[39][16] = 4;
        pixel_data[39][17] = 4;
        pixel_data[39][18] = 4;
        pixel_data[39][19] = 4;
        pixel_data[39][20] = 4;
        pixel_data[39][21] = 4;
        pixel_data[39][22] = 4;
        pixel_data[39][23] = 4;
        pixel_data[39][24] = 4;
        pixel_data[39][25] = 4;
        pixel_data[39][26] = 4;
        pixel_data[39][27] = 4;
        pixel_data[39][28] = 4;
        pixel_data[39][29] = 4;
        pixel_data[39][30] = 4;
        pixel_data[39][31] = 4;
        pixel_data[39][32] = 3;
        pixel_data[39][33] = 3;
        pixel_data[39][34] = 3;
        pixel_data[39][35] = 4;
        pixel_data[39][36] = 4;
        pixel_data[39][37] = 4;
        pixel_data[39][38] = 4;
        pixel_data[39][39] = 4;
        pixel_data[39][40] = 4;
        pixel_data[39][41] = 4;
        pixel_data[39][42] = 4;
        pixel_data[39][43] = 15;
        pixel_data[39][44] = 8;
        pixel_data[39][45] = 8;
        pixel_data[39][46] = 8;
        pixel_data[39][47] = 8;
        pixel_data[39][48] = 8;
        pixel_data[39][49] = 8; // y=39
        pixel_data[40][0] = 0;
        pixel_data[40][1] = 13;
        pixel_data[40][2] = 8;
        pixel_data[40][3] = 8;
        pixel_data[40][4] = 8;
        pixel_data[40][5] = 8;
        pixel_data[40][6] = 8;
        pixel_data[40][7] = 8;
        pixel_data[40][8] = 5;
        pixel_data[40][9] = 4;
        pixel_data[40][10] = 4;
        pixel_data[40][11] = 4;
        pixel_data[40][12] = 4;
        pixel_data[40][13] = 4;
        pixel_data[40][14] = 4;
        pixel_data[40][15] = 4;
        pixel_data[40][16] = 4;
        pixel_data[40][17] = 4;
        pixel_data[40][18] = 4;
        pixel_data[40][19] = 4;
        pixel_data[40][20] = 4;
        pixel_data[40][21] = 4;
        pixel_data[40][22] = 4;
        pixel_data[40][23] = 4;
        pixel_data[40][24] = 4;
        pixel_data[40][25] = 4;
        pixel_data[40][26] = 4;
        pixel_data[40][27] = 4;
        pixel_data[40][28] = 4;
        pixel_data[40][29] = 4;
        pixel_data[40][30] = 4;
        pixel_data[40][31] = 4;
        pixel_data[40][32] = 4;
        pixel_data[40][33] = 4;
        pixel_data[40][34] = 4;
        pixel_data[40][35] = 4;
        pixel_data[40][36] = 4;
        pixel_data[40][37] = 4;
        pixel_data[40][38] = 4;
        pixel_data[40][39] = 4;
        pixel_data[40][40] = 4;
        pixel_data[40][41] = 4;
        pixel_data[40][42] = 5;
        pixel_data[40][43] = 8;
        pixel_data[40][44] = 8;
        pixel_data[40][45] = 8;
        pixel_data[40][46] = 8;
        pixel_data[40][47] = 8;
        pixel_data[40][48] = 8;
        pixel_data[40][49] = 8; // y=40
        pixel_data[41][0] = 0;
        pixel_data[41][1] = 1;
        pixel_data[41][2] = 8;
        pixel_data[41][3] = 8;
        pixel_data[41][4] = 8;
        pixel_data[41][5] = 8;
        pixel_data[41][6] = 8;
        pixel_data[41][7] = 8;
        pixel_data[41][8] = 8;
        pixel_data[41][9] = 5;
        pixel_data[41][10] = 4;
        pixel_data[41][11] = 4;
        pixel_data[41][12] = 4;
        pixel_data[41][13] = 4;
        pixel_data[41][14] = 4;
        pixel_data[41][15] = 4;
        pixel_data[41][16] = 4;
        pixel_data[41][17] = 4;
        pixel_data[41][18] = 4;
        pixel_data[41][19] = 4;
        pixel_data[41][20] = 4;
        pixel_data[41][21] = 4;
        pixel_data[41][22] = 4;
        pixel_data[41][23] = 4;
        pixel_data[41][24] = 4;
        pixel_data[41][25] = 4;
        pixel_data[41][26] = 4;
        pixel_data[41][27] = 4;
        pixel_data[41][28] = 4;
        pixel_data[41][29] = 4;
        pixel_data[41][30] = 4;
        pixel_data[41][31] = 4;
        pixel_data[41][32] = 4;
        pixel_data[41][33] = 4;
        pixel_data[41][34] = 4;
        pixel_data[41][35] = 4;
        pixel_data[41][36] = 4;
        pixel_data[41][37] = 4;
        pixel_data[41][38] = 4;
        pixel_data[41][39] = 4;
        pixel_data[41][40] = 4;
        pixel_data[41][41] = 5;
        pixel_data[41][42] = 8;
        pixel_data[41][43] = 8;
        pixel_data[41][44] = 8;
        pixel_data[41][45] = 8;
        pixel_data[41][46] = 8;
        pixel_data[41][47] = 8;
        pixel_data[41][48] = 8;
        pixel_data[41][49] = 8; // y=41
        pixel_data[42][0] = 0;
        pixel_data[42][1] = 1;
        pixel_data[42][2] = 11;
        pixel_data[42][3] = 8;
        pixel_data[42][4] = 8;
        pixel_data[42][5] = 8;
        pixel_data[42][6] = 8;
        pixel_data[42][7] = 8;
        pixel_data[42][8] = 8;
        pixel_data[42][9] = 8;
        pixel_data[42][10] = 5;
        pixel_data[42][11] = 4;
        pixel_data[42][12] = 3;
        pixel_data[42][13] = 4;
        pixel_data[42][14] = 4;
        pixel_data[42][15] = 4;
        pixel_data[42][16] = 4;
        pixel_data[42][17] = 4;
        pixel_data[42][18] = 4;
        pixel_data[42][19] = 4;
        pixel_data[42][20] = 4;
        pixel_data[42][21] = 4;
        pixel_data[42][22] = 4;
        pixel_data[42][23] = 4;
        pixel_data[42][24] = 4;
        pixel_data[42][25] = 4;
        pixel_data[42][26] = 4;
        pixel_data[42][27] = 4;
        pixel_data[42][28] = 4;
        pixel_data[42][29] = 4;
        pixel_data[42][30] = 4;
        pixel_data[42][31] = 4;
        pixel_data[42][32] = 4;
        pixel_data[42][33] = 4;
        pixel_data[42][34] = 4;
        pixel_data[42][35] = 4;
        pixel_data[42][36] = 4;
        pixel_data[42][37] = 4;
        pixel_data[42][38] = 4;
        pixel_data[42][39] = 4;
        pixel_data[42][40] = 5;
        pixel_data[42][41] = 8;
        pixel_data[42][42] = 8;
        pixel_data[42][43] = 8;
        pixel_data[42][44] = 8;
        pixel_data[42][45] = 8;
        pixel_data[42][46] = 8;
        pixel_data[42][47] = 8;
        pixel_data[42][48] = 8;
        pixel_data[42][49] = 8; // y=42
        pixel_data[43][0] = 0;
        pixel_data[43][1] = 2;
        pixel_data[43][2] = 11;
        pixel_data[43][3] = 8;
        pixel_data[43][4] = 8;
        pixel_data[43][5] = 8;
        pixel_data[43][6] = 8;
        pixel_data[43][7] = 8;
        pixel_data[43][8] = 8;
        pixel_data[43][9] = 8;
        pixel_data[43][10] = 8;
        pixel_data[43][11] = 5;
        pixel_data[43][12] = 6;
        pixel_data[43][13] = 4;
        pixel_data[43][14] = 4;
        pixel_data[43][15] = 4;
        pixel_data[43][16] = 4;
        pixel_data[43][17] = 4;
        pixel_data[43][18] = 4;
        pixel_data[43][19] = 4;
        pixel_data[43][20] = 4;
        pixel_data[43][21] = 4;
        pixel_data[43][22] = 4;
        pixel_data[43][23] = 4;
        pixel_data[43][24] = 4;
        pixel_data[43][25] = 15;
        pixel_data[43][26] = 4;
        pixel_data[43][27] = 4;
        pixel_data[43][28] = 4;
        pixel_data[43][29] = 4;
        pixel_data[43][30] = 4;
        pixel_data[43][31] = 4;
        pixel_data[43][32] = 4;
        pixel_data[43][33] = 4;
        pixel_data[43][34] = 4;
        pixel_data[43][35] = 4;
        pixel_data[43][36] = 4;
        pixel_data[43][37] = 4;
        pixel_data[43][38] = 3;
        pixel_data[43][39] = 5;
        pixel_data[43][40] = 8;
        pixel_data[43][41] = 8;
        pixel_data[43][42] = 8;
        pixel_data[43][43] = 8;
        pixel_data[43][44] = 8;
        pixel_data[43][45] = 8;
        pixel_data[43][46] = 8;
        pixel_data[43][47] = 8;
        pixel_data[43][48] = 8;
        pixel_data[43][49] = 11; // y=43
        pixel_data[44][0] = 1;
        pixel_data[44][1] = 2;
        pixel_data[44][2] = 11;
        pixel_data[44][3] = 8;
        pixel_data[44][4] = 8;
        pixel_data[44][5] = 8;
        pixel_data[44][6] = 8;
        pixel_data[44][7] = 8;
        pixel_data[44][8] = 8;
        pixel_data[44][9] = 8;
        pixel_data[44][10] = 8;
        pixel_data[44][11] = 8;
        pixel_data[44][12] = 11;
        pixel_data[44][13] = 6;
        pixel_data[44][14] = 3;
        pixel_data[44][15] = 4;
        pixel_data[44][16] = 4;
        pixel_data[44][17] = 4;
        pixel_data[44][18] = 4;
        pixel_data[44][19] = 4;
        pixel_data[44][20] = 4;
        pixel_data[44][21] = 4;
        pixel_data[44][22] = 4;
        pixel_data[44][23] = 3;
        pixel_data[44][24] = 4;
        pixel_data[44][25] = 9;
        pixel_data[44][26] = 4;
        pixel_data[44][27] = 3;
        pixel_data[44][28] = 4;
        pixel_data[44][29] = 4;
        pixel_data[44][30] = 4;
        pixel_data[44][31] = 4;
        pixel_data[44][32] = 4;
        pixel_data[44][33] = 4;
        pixel_data[44][34] = 4;
        pixel_data[44][35] = 3;
        pixel_data[44][36] = 3;
        pixel_data[44][37] = 6;
        pixel_data[44][38] = 8;
        pixel_data[44][39] = 8;
        pixel_data[44][40] = 8;
        pixel_data[44][41] = 8;
        pixel_data[44][42] = 8;
        pixel_data[44][43] = 8;
        pixel_data[44][44] = 8;
        pixel_data[44][45] = 8;
        pixel_data[44][46] = 8;
        pixel_data[44][47] = 8;
        pixel_data[44][48] = 8;
        pixel_data[44][49] = 1; // y=44
        pixel_data[45][0] = 13;
        pixel_data[45][1] = 0;
        pixel_data[45][2] = 13;
        pixel_data[45][3] = 8;
        pixel_data[45][4] = 8;
        pixel_data[45][5] = 8;
        pixel_data[45][6] = 8;
        pixel_data[45][7] = 8;
        pixel_data[45][8] = 8;
        pixel_data[45][9] = 8;
        pixel_data[45][10] = 8;
        pixel_data[45][11] = 11;
        pixel_data[45][12] = 2;
        pixel_data[45][13] = 8;
        pixel_data[45][14] = 5;
        pixel_data[45][15] = 4;
        pixel_data[45][16] = 4;
        pixel_data[45][17] = 4;
        pixel_data[45][18] = 4;
        pixel_data[45][19] = 4;
        pixel_data[45][20] = 4;
        pixel_data[45][21] = 4;
        pixel_data[45][22] = 4;
        pixel_data[45][23] = 15;
        pixel_data[45][24] = 9;
        pixel_data[45][25] = 10;
        pixel_data[45][26] = 9;
        pixel_data[45][27] = 15;
        pixel_data[45][28] = 4;
        pixel_data[45][29] = 4;
        pixel_data[45][30] = 4;
        pixel_data[45][31] = 4;
        pixel_data[45][32] = 4;
        pixel_data[45][33] = 4;
        pixel_data[45][34] = 15;
        pixel_data[45][35] = 9;
        pixel_data[45][36] = 11;
        pixel_data[45][37] = 8;
        pixel_data[45][38] = 8;
        pixel_data[45][39] = 8;
        pixel_data[45][40] = 8;
        pixel_data[45][41] = 8;
        pixel_data[45][42] = 8;
        pixel_data[45][43] = 8;
        pixel_data[45][44] = 8;
        pixel_data[45][45] = 8;
        pixel_data[45][46] = 8;
        pixel_data[45][47] = 8;
        pixel_data[45][48] = 13;
        pixel_data[45][49] = 2; // y=45
        pixel_data[46][0] = 2;
        pixel_data[46][1] = 2;
        pixel_data[46][2] = 2;
        pixel_data[46][3] = 13;
        pixel_data[46][4] = 8;
        pixel_data[46][5] = 8;
        pixel_data[46][6] = 8;
        pixel_data[46][7] = 8;
        pixel_data[46][8] = 8;
        pixel_data[46][9] = 8;
        pixel_data[46][10] = 8;
        pixel_data[46][11] = 1;
        pixel_data[46][12] = 0;
        pixel_data[46][13] = 13;
        pixel_data[46][14] = 8;
        pixel_data[46][15] = 8;
        pixel_data[46][16] = 5;
        pixel_data[46][17] = 4;
        pixel_data[46][18] = 4;
        pixel_data[46][19] = 4;
        pixel_data[46][20] = 4;
        pixel_data[46][21] = 4;
        pixel_data[46][22] = 4;
        pixel_data[46][23] = 4;
        pixel_data[46][24] = 9;
        pixel_data[46][25] = 14;
        pixel_data[46][26] = 10;
        pixel_data[46][27] = 4;
        pixel_data[46][28] = 3;
        pixel_data[46][29] = 4;
        pixel_data[46][30] = 4;
        pixel_data[46][31] = 4;
        pixel_data[46][32] = 6;
        pixel_data[46][33] = 3;
        pixel_data[46][34] = 5;
        pixel_data[46][35] = 13;
        pixel_data[46][36] = 1;
        pixel_data[46][37] = 8;
        pixel_data[46][38] = 8;
        pixel_data[46][39] = 8;
        pixel_data[46][40] = 8;
        pixel_data[46][41] = 8;
        pixel_data[46][42] = 8;
        pixel_data[46][43] = 8;
        pixel_data[46][44] = 8;
        pixel_data[46][45] = 8;
        pixel_data[46][46] = 11;
        pixel_data[46][47] = 1;
        pixel_data[46][48] = 2;
        pixel_data[46][49] = 1; // y=46
        pixel_data[47][0] = 0;
        pixel_data[47][1] = 11;
        pixel_data[47][2] = 0;
        pixel_data[47][3] = 1;
        pixel_data[47][4] = 11;
        pixel_data[47][5] = 15;
        pixel_data[47][6] = 8;
        pixel_data[47][7] = 8;
        pixel_data[47][8] = 8;
        pixel_data[47][9] = 8;
        pixel_data[47][10] = 13;
        pixel_data[47][11] = 2;
        pixel_data[47][12] = 0;
        pixel_data[47][13] = 1;
        pixel_data[47][14] = 11;
        pixel_data[47][15] = 15;
        pixel_data[47][16] = 8;
        pixel_data[47][17] = 8;
        pixel_data[47][18] = 5;
        pixel_data[47][19] = 5;
        pixel_data[47][20] = 4;
        pixel_data[47][21] = 4;
        pixel_data[47][22] = 15;
        pixel_data[47][23] = 9;
        pixel_data[47][24] = 9;
        pixel_data[47][25] = 14;
        pixel_data[47][26] = 15;
        pixel_data[47][27] = 10;
        pixel_data[47][28] = 3;
        pixel_data[47][29] = 15;
        pixel_data[47][30] = 15;
        pixel_data[47][31] = 5;
        pixel_data[47][32] = 15;
        pixel_data[47][33] = 8;
        pixel_data[47][34] = 11;
        pixel_data[47][35] = 2;
        pixel_data[47][36] = 2;
        pixel_data[47][37] = 13;
        pixel_data[47][38] = 8;
        pixel_data[47][39] = 15;
        pixel_data[47][40] = 8;
        pixel_data[47][41] = 15;
        pixel_data[47][42] = 15;
        pixel_data[47][43] = 15;
        pixel_data[47][44] = 8;
        pixel_data[47][45] = 13;
        pixel_data[47][46] = 2;
        pixel_data[47][47] = 0;
        pixel_data[47][48] = 0;
        pixel_data[47][49] = 2; // y=47
        pixel_data[48][0] = 0;
        pixel_data[48][1] = 0;
        pixel_data[48][2] = 5;
        pixel_data[48][3] = 0;
        pixel_data[48][4] = 13;
        pixel_data[48][5] = 11;
        pixel_data[48][6] = 11;
        pixel_data[48][7] = 11;
        pixel_data[48][8] = 11;
        pixel_data[48][9] = 11;
        pixel_data[48][10] = 1;
        pixel_data[48][11] = 0;
        pixel_data[48][12] = 1;
        pixel_data[48][13] = 2;
        pixel_data[48][14] = 13;
        pixel_data[48][15] = 11;
        pixel_data[48][16] = 8;
        pixel_data[48][17] = 8;
        pixel_data[48][18] = 8;
        pixel_data[48][19] = 8;
        pixel_data[48][20] = 8;
        pixel_data[48][21] = 15;
        pixel_data[48][22] = 11;
        pixel_data[48][23] = 10;
        pixel_data[48][24] = 14;
        pixel_data[48][25] = 14;
        pixel_data[48][26] = 14;
        pixel_data[48][27] = 10;
        pixel_data[48][28] = 9;
        pixel_data[48][29] = 11;
        pixel_data[48][30] = 11;
        pixel_data[48][31] = 11;
        pixel_data[48][32] = 11;
        pixel_data[48][33] = 11;
        pixel_data[48][34] = 1;
        pixel_data[48][35] = 0;
        pixel_data[48][36] = 0;
        pixel_data[48][37] = 1;
        pixel_data[48][38] = 8;
        pixel_data[48][39] = 11;
        pixel_data[48][40] = 11;
        pixel_data[48][41] = 11;
        pixel_data[48][42] = 11;
        pixel_data[48][43] = 8;
        pixel_data[48][44] = 11;
        pixel_data[48][45] = 2;
        pixel_data[48][46] = 0;
        pixel_data[48][47] = 11;
        pixel_data[48][48] = 0;
        pixel_data[48][49] = 0; // y=48
        pixel_data[49][0] = 0;
        pixel_data[49][1] = 0;
        pixel_data[49][2] = 0;
        pixel_data[49][3] = 1;
        pixel_data[49][4] = 0;
        pixel_data[49][5] = 2;
        pixel_data[49][6] = 1;
        pixel_data[49][7] = 13;
        pixel_data[49][8] = 1;
        pixel_data[49][9] = 2;
        pixel_data[49][10] = 0;
        pixel_data[49][11] = 2;
        pixel_data[49][12] = 0;
        pixel_data[49][13] = 1;
        pixel_data[49][14] = 0;
        pixel_data[49][15] = 2;
        pixel_data[49][16] = 11;
        pixel_data[49][17] = 13;
        pixel_data[49][18] = 13;
        pixel_data[49][19] = 11;
        pixel_data[49][20] = 11;
        pixel_data[49][21] = 13;
        pixel_data[49][22] = 1;
        pixel_data[49][23] = 0;
        pixel_data[49][24] = 0;
        pixel_data[49][25] = 0;
        pixel_data[49][26] = 0;
        pixel_data[49][27] = 0;
        pixel_data[49][28] = 0;
        pixel_data[49][29] = 2;
        pixel_data[49][30] = 2;
        pixel_data[49][31] = 1;
        pixel_data[49][32] = 2;
        pixel_data[49][33] = 0;
        pixel_data[49][34] = 0;
        pixel_data[49][35] = 2;
        pixel_data[49][36] = 0;
        pixel_data[49][37] = 0;
        pixel_data[49][38] = 0;
        pixel_data[49][39] = 2;
        pixel_data[49][40] = 2;
        pixel_data[49][41] = 2;
        pixel_data[49][42] = 2;
        pixel_data[49][43] = 0;
        pixel_data[49][44] = 0;
        pixel_data[49][45] = 0;
        pixel_data[49][46] = 2;
        pixel_data[49][47] = 0;
        pixel_data[49][48] = 0;
        pixel_data[49][49] = 0; // y=49
    end
endmodule